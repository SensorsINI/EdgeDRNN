module edgedrnn_wrapper #(
    parameter integer C_S_AXI_DATA_WIDTH = 32,
    parameter integer C_S_AXI_ADDR_WIDTH = 7,
    parameter integer NUM_PE             = 8, // >= 2
    parameter integer ACT_INT_BW         = 8,
    parameter integer ACT_FRA_BW         = 8,
    parameter integer W_INT_BW           = 1,
    parameter integer W_FRA_BW           = 7,
    parameter integer NUM_LAYER_BW       = 2,
    parameter integer LAYER_SIZE_BW      = 10,  
    parameter integer DTH_BW             = 10,
    parameter integer NZI_BW             = 16,
    parameter integer NZL_FIFO_DEPTH     = 32
    )(
    input  wire                                        clk,
    input  wire                                        rst_n,
    input  wire [C_S_AXI_ADDR_WIDTH-1:0]               s_axi_awaddr,
    input  wire [2:0]                                  s_axi_awprot,
    input  wire                                        s_axi_awvalid,
    output wire                                        s_axi_awready,
    input  wire [C_S_AXI_DATA_WIDTH-1:0]               s_axi_wdata,
    input  wire [(C_S_AXI_DATA_WIDTH/8)-1:0]           s_axi_wstrb,
    input  wire                                        s_axi_wvalid,
    output wire                                        s_axi_wready,
    output wire [1:0]                                  s_axi_bresp,
    output wire                                        s_axi_bvalid,
    input  wire                                        s_axi_bready,
    input  wire [C_S_AXI_ADDR_WIDTH-1:0]               s_axi_araddr,
    input  wire [2:0]                                  s_axi_arprot,
    input  wire                                        s_axi_arvalid,
    output wire                                        s_axi_arready,
    output wire [C_S_AXI_DATA_WIDTH-1:0]               s_axi_rdata,
    output wire [1:0]                                  s_axi_rresp,
    output wire                                        s_axi_rvalid,
    input  wire                                        s_axi_rready,
    input  wire                                        s_inp_axis_tvalid,
    output wire                                        s_inp_axis_tready,
    input  wire [NUM_PE*(ACT_INT_BW + ACT_FRA_BW)-1:0] s_inp_axis_tdata,
    input  wire                                        s_inp_axis_tlast,
    input  wire                                        s_w_axis_tvalid,
    output wire                                        s_w_axis_tready,
    input  wire [NUM_PE*(W_INT_BW + W_FRA_BW)-1:0]     s_w_axis_tdata,
    input  wire                                        s_w_axis_tlast,
    output wire                                        m_inst_axis_tvalid,
    input  wire                                        m_inst_axis_tready,
    output wire [80-1:0]                               m_inst_axis_tdata,
    output wire                                        m_inst_axis_tlast,
    output wire                                        m_out_axis_tvalid,
    input  wire                                        m_out_axis_tready,
    output wire [NUM_PE*(ACT_INT_BW + ACT_FRA_BW)-1:0] m_out_axis_tdata,
    output wire                                        m_out_axis_tlast
    );
    
    edgedrnn # (
        .C_S_AXI_DATA_WIDTH (C_S_AXI_DATA_WIDTH),
        .C_S_AXI_ADDR_WIDTH (C_S_AXI_ADDR_WIDTH),
        .NUM_PE             (NUM_PE            ),
        .ACT_INT_BW         (ACT_INT_BW        ),
        .ACT_FRA_BW         (ACT_FRA_BW        ),
        .W_INT_BW           (W_INT_BW          ),
        .W_FRA_BW           (W_FRA_BW          ),
        .NUM_LAYER_BW       (NUM_LAYER_BW      ),
        .LAYER_SIZE_BW      (LAYER_SIZE_BW     ),
        .DTH_BW             (DTH_BW            ),
        .NZI_BW             (NZI_BW            ),
        .NZL_FIFO_DEPTH     (NZL_FIFO_DEPTH    )     
    ) i_edgedrnn (
        .clk                (clk               ),
        .rst_n              (rst_n             ),
        .s_axi_awaddr       (s_axi_awaddr      ),
        .s_axi_awprot       (s_axi_awprot      ),
        .s_axi_awvalid      (s_axi_awvalid     ),
        .s_axi_awready      (s_axi_awready     ),
        .s_axi_wdata        (s_axi_wdata       ),
        .s_axi_wstrb        (s_axi_wstrb       ),
        .s_axi_wvalid       (s_axi_wvalid      ),
        .s_axi_wready       (s_axi_wready      ),
        .s_axi_bresp        (s_axi_bresp       ),
        .s_axi_bvalid       (s_axi_bvalid      ),
        .s_axi_bready       (s_axi_bready      ),
        .s_axi_araddr       (s_axi_araddr      ),
        .s_axi_arprot       (s_axi_arprot      ),
        .s_axi_arvalid      (s_axi_arvalid     ),
        .s_axi_arready      (s_axi_arready     ),
        .s_axi_rdata        (s_axi_rdata       ),
        .s_axi_rresp        (s_axi_rresp       ),
        .s_axi_rvalid       (s_axi_rvalid      ),
        .s_axi_rready       (s_axi_rready      ),
        .s_inp_axis_tvalid  (s_inp_axis_tvalid ),
        .s_inp_axis_tready  (s_inp_axis_tready ),
        .s_inp_axis_tdata   (s_inp_axis_tdata  ),
        .s_inp_axis_tlast   (s_inp_axis_tlast  ),  
        .s_w_axis_tvalid    (s_w_axis_tvalid   ),
        .s_w_axis_tready    (s_w_axis_tready   ),
        .s_w_axis_tdata     (s_w_axis_tdata    ),
        .s_w_axis_tlast     (s_w_axis_tlast    ),  
        .m_inst_axis_tvalid (m_inst_axis_tvalid),
        .m_inst_axis_tready (m_inst_axis_tready),
        .m_inst_axis_tdata  (m_inst_axis_tdata ),
        .m_inst_axis_tlast  (m_inst_axis_tlast ),
        .m_out_axis_tvalid  (m_out_axis_tvalid ),
        .m_out_axis_tready  (m_out_axis_tready ),
        .m_out_axis_tdata   (m_out_axis_tdata  ),
        .m_out_axis_tlast   (m_out_axis_tlast  )
    );

    endmodule
