module tanh_lut #(
   NUM_PE     = 1,
   ACT_INT_BW = 8,
   ACT_FRA_BW = 8
   )(
   input  logic signed [NUM_PE-1:0][ACT_INT_BW+ACT_FRA_BW-1:0] in,
   output logic signed [NUM_PE-1:0][ACT_INT_BW+ACT_FRA_BW-1:0] out
   );
   
   localparam ACT_BW = ACT_INT_BW + ACT_FRA_BW;
   logic signed [NUM_PE-1:0][ACT_BW-1:0] lut_in;
   logic signed [NUM_PE-1:0][ACT_BW-1:0] lut_out;
   
   assign out = lut_out;

   always_comb begin
      for (int unsigned i = 0; i < NUM_PE; i = i + 1) begin
         lut_out[i] = '0;
         lut_in[i] = in[i];
         if ($signed(in[i]) > $signed(530)) begin // 2047
            lut_out[i] = $signed(256);
         end else if ($signed(in[i]) < $signed(-530)) begin //-2048
            lut_out[i] = $signed(-256);
         end else begin
            case($signed(lut_in[i]))
               -530 : lut_out[i] = -240;
               -529 : lut_out[i] = -240;
               -528 : lut_out[i] = -240;
               -527 : lut_out[i] = -240;
               -526 : lut_out[i] = -240;
               -525 : lut_out[i] = -240;
               -524 : lut_out[i] = -240;
               -523 : lut_out[i] = -240;
               -522 : lut_out[i] = -240;
               -521 : lut_out[i] = -240;
               -520 : lut_out[i] = -240;
               -519 : lut_out[i] = -240;
               -518 : lut_out[i] = -240;
               -517 : lut_out[i] = -240;
               -516 : lut_out[i] = -240;
               -515 : lut_out[i] = -240;
               -514 : lut_out[i] = -240;
               -513 : lut_out[i] = -240;
               -512 : lut_out[i] = -240;
               -511 : lut_out[i] = -240;
               -510 : lut_out[i] = -240;
               -509 : lut_out[i] = -240;
               -508 : lut_out[i] = -240;
               -507 : lut_out[i] = -240;
               -506 : lut_out[i] = -240;
               -505 : lut_out[i] = -240;
               -504 : lut_out[i] = -240;
               -503 : lut_out[i] = -240;
               -502 : lut_out[i] = -240;
               -501 : lut_out[i] = -240;
               -500 : lut_out[i] = -240;
               -499 : lut_out[i] = -240;
               -498 : lut_out[i] = -240;
               -497 : lut_out[i] = -240;
               -496 : lut_out[i] = -240;
               -495 : lut_out[i] = -240;
               -494 : lut_out[i] = -240;
               -493 : lut_out[i] = -240;
               -492 : lut_out[i] = -240;
               -491 : lut_out[i] = -240;
               -490 : lut_out[i] = -240;
               -489 : lut_out[i] = -240;
               -488 : lut_out[i] = -240;
               -487 : lut_out[i] = -240;
               -486 : lut_out[i] = -240;
               -485 : lut_out[i] = -240;
               -484 : lut_out[i] = -240;
               -483 : lut_out[i] = -240;
               -482 : lut_out[i] = -240;
               -481 : lut_out[i] = -240;
               -480 : lut_out[i] = -240;
               -479 : lut_out[i] = -240;
               -478 : lut_out[i] = -240;
               -477 : lut_out[i] = -240;
               -476 : lut_out[i] = -240;
               -475 : lut_out[i] = -240;
               -474 : lut_out[i] = -240;
               -473 : lut_out[i] = -240;
               -472 : lut_out[i] = -240;
               -471 : lut_out[i] = -240;
               -470 : lut_out[i] = -240;
               -469 : lut_out[i] = -240;
               -468 : lut_out[i] = -240;
               -467 : lut_out[i] = -240;
               -466 : lut_out[i] = -240;
               -465 : lut_out[i] = -240;
               -464 : lut_out[i] = -240;
               -463 : lut_out[i] = -240;
               -462 : lut_out[i] = -240;
               -461 : lut_out[i] = -240;
               -460 : lut_out[i] = -240;
               -459 : lut_out[i] = -240;
               -458 : lut_out[i] = -240;
               -457 : lut_out[i] = -240;
               -456 : lut_out[i] = -240;
               -455 : lut_out[i] = -240;
               -454 : lut_out[i] = -240;
               -453 : lut_out[i] = -240;
               -452 : lut_out[i] = -240;
               -451 : lut_out[i] = -240;
               -450 : lut_out[i] = -240;
               -449 : lut_out[i] = -240;
               -448 : lut_out[i] = -240;
               -447 : lut_out[i] = -240;
               -446 : lut_out[i] = -240;
               -445 : lut_out[i] = -240;
               -444 : lut_out[i] = -240;
               -443 : lut_out[i] = -240;
               -442 : lut_out[i] = -240;
               -441 : lut_out[i] = -240;
               -440 : lut_out[i] = -240;
               -439 : lut_out[i] = -240;
               -438 : lut_out[i] = -240;
               -437 : lut_out[i] = -240;
               -436 : lut_out[i] = -240;
               -435 : lut_out[i] = -240;
               -434 : lut_out[i] = -240;
               -433 : lut_out[i] = -240;
               -432 : lut_out[i] = -240;
               -431 : lut_out[i] = -240;
               -430 : lut_out[i] = -240;
               -429 : lut_out[i] = -240;
               -428 : lut_out[i] = -240;
               -427 : lut_out[i] = -240;
               -426 : lut_out[i] = -240;
               -425 : lut_out[i] = -240;
               -424 : lut_out[i] = -240;
               -423 : lut_out[i] = -240;
               -422 : lut_out[i] = -240;
               -421 : lut_out[i] = -240;
               -420 : lut_out[i] = -240;
               -419 : lut_out[i] = -240;
               -418 : lut_out[i] = -240;
               -417 : lut_out[i] = -240;
               -416 : lut_out[i] = -240;
               -415 : lut_out[i] = -240;
               -414 : lut_out[i] = -240;
               -413 : lut_out[i] = -240;
               -412 : lut_out[i] = -240;
               -411 : lut_out[i] = -240;
               -410 : lut_out[i] = -240;
               -409 : lut_out[i] = -240;
               -408 : lut_out[i] = -240;
               -407 : lut_out[i] = -240;
               -406 : lut_out[i] = -240;
               -405 : lut_out[i] = -240;
               -404 : lut_out[i] = -240;
               -403 : lut_out[i] = -240;
               -402 : lut_out[i] = -240;
               -401 : lut_out[i] = -240;
               -400 : lut_out[i] = -240;
               -399 : lut_out[i] = -240;
               -398 : lut_out[i] = -240;
               -397 : lut_out[i] = -240;
               -396 : lut_out[i] = -240;
               -395 : lut_out[i] = -240;
               -394 : lut_out[i] = -240;
               -393 : lut_out[i] = -240;
               -392 : lut_out[i] = -240;
               -391 : lut_out[i] = -240;
               -390 : lut_out[i] = -240;
               -389 : lut_out[i] = -240;
               -388 : lut_out[i] = -240;
               -387 : lut_out[i] = -240;
               -386 : lut_out[i] = -240;
               -385 : lut_out[i] = -224;
               -384 : lut_out[i] = -224;
               -383 : lut_out[i] = -224;
               -382 : lut_out[i] = -224;
               -381 : lut_out[i] = -224;
               -380 : lut_out[i] = -224;
               -379 : lut_out[i] = -224;
               -378 : lut_out[i] = -224;
               -377 : lut_out[i] = -224;
               -376 : lut_out[i] = -224;
               -375 : lut_out[i] = -224;
               -374 : lut_out[i] = -224;
               -373 : lut_out[i] = -224;
               -372 : lut_out[i] = -224;
               -371 : lut_out[i] = -224;
               -370 : lut_out[i] = -224;
               -369 : lut_out[i] = -224;
               -368 : lut_out[i] = -224;
               -367 : lut_out[i] = -224;
               -366 : lut_out[i] = -224;
               -365 : lut_out[i] = -224;
               -364 : lut_out[i] = -224;
               -363 : lut_out[i] = -224;
               -362 : lut_out[i] = -224;
               -361 : lut_out[i] = -224;
               -360 : lut_out[i] = -224;
               -359 : lut_out[i] = -224;
               -358 : lut_out[i] = -224;
               -357 : lut_out[i] = -224;
               -356 : lut_out[i] = -224;
               -355 : lut_out[i] = -224;
               -354 : lut_out[i] = -224;
               -353 : lut_out[i] = -224;
               -352 : lut_out[i] = -224;
               -351 : lut_out[i] = -224;
               -350 : lut_out[i] = -224;
               -349 : lut_out[i] = -224;
               -348 : lut_out[i] = -224;
               -347 : lut_out[i] = -224;
               -346 : lut_out[i] = -224;
               -345 : lut_out[i] = -224;
               -344 : lut_out[i] = -224;
               -343 : lut_out[i] = -224;
               -342 : lut_out[i] = -224;
               -341 : lut_out[i] = -224;
               -340 : lut_out[i] = -224;
               -339 : lut_out[i] = -224;
               -338 : lut_out[i] = -224;
               -337 : lut_out[i] = -224;
               -336 : lut_out[i] = -224;
               -335 : lut_out[i] = -224;
               -334 : lut_out[i] = -224;
               -333 : lut_out[i] = -224;
               -332 : lut_out[i] = -224;
               -331 : lut_out[i] = -224;
               -330 : lut_out[i] = -224;
               -329 : lut_out[i] = -224;
               -328 : lut_out[i] = -224;
               -327 : lut_out[i] = -224;
               -326 : lut_out[i] = -224;
               -325 : lut_out[i] = -224;
               -324 : lut_out[i] = -224;
               -323 : lut_out[i] = -224;
               -322 : lut_out[i] = -224;
               -321 : lut_out[i] = -224;
               -320 : lut_out[i] = -224;
               -319 : lut_out[i] = -224;
               -318 : lut_out[i] = -224;
               -317 : lut_out[i] = -224;
               -316 : lut_out[i] = -224;
               -315 : lut_out[i] = -208;
               -314 : lut_out[i] = -208;
               -313 : lut_out[i] = -208;
               -312 : lut_out[i] = -208;
               -311 : lut_out[i] = -208;
               -310 : lut_out[i] = -208;
               -309 : lut_out[i] = -208;
               -308 : lut_out[i] = -208;
               -307 : lut_out[i] = -208;
               -306 : lut_out[i] = -208;
               -305 : lut_out[i] = -208;
               -304 : lut_out[i] = -208;
               -303 : lut_out[i] = -208;
               -302 : lut_out[i] = -208;
               -301 : lut_out[i] = -208;
               -300 : lut_out[i] = -208;
               -299 : lut_out[i] = -208;
               -298 : lut_out[i] = -208;
               -297 : lut_out[i] = -208;
               -296 : lut_out[i] = -208;
               -295 : lut_out[i] = -208;
               -294 : lut_out[i] = -208;
               -293 : lut_out[i] = -208;
               -292 : lut_out[i] = -208;
               -291 : lut_out[i] = -208;
               -290 : lut_out[i] = -208;
               -289 : lut_out[i] = -208;
               -288 : lut_out[i] = -208;
               -287 : lut_out[i] = -208;
               -286 : lut_out[i] = -208;
               -285 : lut_out[i] = -208;
               -284 : lut_out[i] = -208;
               -283 : lut_out[i] = -208;
               -282 : lut_out[i] = -208;
               -281 : lut_out[i] = -208;
               -280 : lut_out[i] = -208;
               -279 : lut_out[i] = -208;
               -278 : lut_out[i] = -208;
               -277 : lut_out[i] = -208;
               -276 : lut_out[i] = -208;
               -275 : lut_out[i] = -208;
               -274 : lut_out[i] = -208;
               -273 : lut_out[i] = -208;
               -272 : lut_out[i] = -208;
               -271 : lut_out[i] = -208;
               -270 : lut_out[i] = -208;
               -269 : lut_out[i] = -208;
               -268 : lut_out[i] = -192;
               -267 : lut_out[i] = -192;
               -266 : lut_out[i] = -192;
               -265 : lut_out[i] = -192;
               -264 : lut_out[i] = -192;
               -263 : lut_out[i] = -192;
               -262 : lut_out[i] = -192;
               -261 : lut_out[i] = -192;
               -260 : lut_out[i] = -192;
               -259 : lut_out[i] = -192;
               -258 : lut_out[i] = -192;
               -257 : lut_out[i] = -192;
               -256 : lut_out[i] = -192;
               -255 : lut_out[i] = -192;
               -254 : lut_out[i] = -192;
               -253 : lut_out[i] = -192;
               -252 : lut_out[i] = -192;
               -251 : lut_out[i] = -192;
               -250 : lut_out[i] = -192;
               -249 : lut_out[i] = -192;
               -248 : lut_out[i] = -192;
               -247 : lut_out[i] = -192;
               -246 : lut_out[i] = -192;
               -245 : lut_out[i] = -192;
               -244 : lut_out[i] = -192;
               -243 : lut_out[i] = -192;
               -242 : lut_out[i] = -192;
               -241 : lut_out[i] = -192;
               -240 : lut_out[i] = -192;
               -239 : lut_out[i] = -192;
               -238 : lut_out[i] = -192;
               -237 : lut_out[i] = -192;
               -236 : lut_out[i] = -192;
               -235 : lut_out[i] = -192;
               -234 : lut_out[i] = -192;
               -233 : lut_out[i] = -192;
               -232 : lut_out[i] = -192;
               -231 : lut_out[i] = -176;
               -230 : lut_out[i] = -176;
               -229 : lut_out[i] = -176;
               -228 : lut_out[i] = -176;
               -227 : lut_out[i] = -176;
               -226 : lut_out[i] = -176;
               -225 : lut_out[i] = -176;
               -224 : lut_out[i] = -176;
               -223 : lut_out[i] = -176;
               -222 : lut_out[i] = -176;
               -221 : lut_out[i] = -176;
               -220 : lut_out[i] = -176;
               -219 : lut_out[i] = -176;
               -218 : lut_out[i] = -176;
               -217 : lut_out[i] = -176;
               -216 : lut_out[i] = -176;
               -215 : lut_out[i] = -176;
               -214 : lut_out[i] = -176;
               -213 : lut_out[i] = -176;
               -212 : lut_out[i] = -176;
               -211 : lut_out[i] = -176;
               -210 : lut_out[i] = -176;
               -209 : lut_out[i] = -176;
               -208 : lut_out[i] = -176;
               -207 : lut_out[i] = -176;
               -206 : lut_out[i] = -176;
               -205 : lut_out[i] = -176;
               -204 : lut_out[i] = -176;
               -203 : lut_out[i] = -176;
               -202 : lut_out[i] = -176;
               -201 : lut_out[i] = -160;
               -200 : lut_out[i] = -160;
               -199 : lut_out[i] = -160;
               -198 : lut_out[i] = -160;
               -197 : lut_out[i] = -160;
               -196 : lut_out[i] = -160;
               -195 : lut_out[i] = -160;
               -194 : lut_out[i] = -160;
               -193 : lut_out[i] = -160;
               -192 : lut_out[i] = -160;
               -191 : lut_out[i] = -160;
               -190 : lut_out[i] = -160;
               -189 : lut_out[i] = -160;
               -188 : lut_out[i] = -160;
               -187 : lut_out[i] = -160;
               -186 : lut_out[i] = -160;
               -185 : lut_out[i] = -160;
               -184 : lut_out[i] = -160;
               -183 : lut_out[i] = -160;
               -182 : lut_out[i] = -160;
               -181 : lut_out[i] = -160;
               -180 : lut_out[i] = -160;
               -179 : lut_out[i] = -160;
               -178 : lut_out[i] = -160;
               -177 : lut_out[i] = -160;
               -176 : lut_out[i] = -160;
               -175 : lut_out[i] = -160;
               -174 : lut_out[i] = -144;
               -173 : lut_out[i] = -144;
               -172 : lut_out[i] = -144;
               -171 : lut_out[i] = -144;
               -170 : lut_out[i] = -144;
               -169 : lut_out[i] = -144;
               -168 : lut_out[i] = -144;
               -167 : lut_out[i] = -144;
               -166 : lut_out[i] = -144;
               -165 : lut_out[i] = -144;
               -164 : lut_out[i] = -144;
               -163 : lut_out[i] = -144;
               -162 : lut_out[i] = -144;
               -161 : lut_out[i] = -144;
               -160 : lut_out[i] = -144;
               -159 : lut_out[i] = -144;
               -158 : lut_out[i] = -144;
               -157 : lut_out[i] = -144;
               -156 : lut_out[i] = -144;
               -155 : lut_out[i] = -144;
               -154 : lut_out[i] = -144;
               -153 : lut_out[i] = -144;
               -152 : lut_out[i] = -144;
               -151 : lut_out[i] = -128;
               -150 : lut_out[i] = -128;
               -149 : lut_out[i] = -128;
               -148 : lut_out[i] = -128;
               -147 : lut_out[i] = -128;
               -146 : lut_out[i] = -128;
               -145 : lut_out[i] = -128;
               -144 : lut_out[i] = -128;
               -143 : lut_out[i] = -128;
               -142 : lut_out[i] = -128;
               -141 : lut_out[i] = -128;
               -140 : lut_out[i] = -128;
               -139 : lut_out[i] = -128;
               -138 : lut_out[i] = -128;
               -137 : lut_out[i] = -128;
               -136 : lut_out[i] = -128;
               -135 : lut_out[i] = -128;
               -134 : lut_out[i] = -128;
               -133 : lut_out[i] = -128;
               -132 : lut_out[i] = -128;
               -131 : lut_out[i] = -128;
               -130 : lut_out[i] = -112;
               -129 : lut_out[i] = -112;
               -128 : lut_out[i] = -112;
               -127 : lut_out[i] = -112;
               -126 : lut_out[i] = -112;
               -125 : lut_out[i] = -112;
               -124 : lut_out[i] = -112;
               -123 : lut_out[i] = -112;
               -122 : lut_out[i] = -112;
               -121 : lut_out[i] = -112;
               -120 : lut_out[i] = -112;
               -119 : lut_out[i] = -112;
               -118 : lut_out[i] = -112;
               -117 : lut_out[i] = -112;
               -116 : lut_out[i] = -112;
               -115 : lut_out[i] = -112;
               -114 : lut_out[i] = -112;
               -113 : lut_out[i] = -112;
               -112 : lut_out[i] = -112;
               -111 : lut_out[i] = -112;
               -110 : lut_out[i] = -96;
               -109 : lut_out[i] = -96;
               -108 : lut_out[i] = -96;
               -107 : lut_out[i] = -96;
               -106 : lut_out[i] = -96;
               -105 : lut_out[i] = -96;
               -104 : lut_out[i] = -96;
               -103 : lut_out[i] = -96;
               -102 : lut_out[i] = -96;
               -101 : lut_out[i] = -96;
               -100 : lut_out[i] = -96;
               -99 : lut_out[i] = -96;
               -98 : lut_out[i] = -96;
               -97 : lut_out[i] = -96;
               -96 : lut_out[i] = -96;
               -95 : lut_out[i] = -96;
               -94 : lut_out[i] = -96;
               -93 : lut_out[i] = -96;
               -92 : lut_out[i] = -96;
               -91 : lut_out[i] = -80;
               -90 : lut_out[i] = -80;
               -89 : lut_out[i] = -80;
               -88 : lut_out[i] = -80;
               -87 : lut_out[i] = -80;
               -86 : lut_out[i] = -80;
               -85 : lut_out[i] = -80;
               -84 : lut_out[i] = -80;
               -83 : lut_out[i] = -80;
               -82 : lut_out[i] = -80;
               -81 : lut_out[i] = -80;
               -80 : lut_out[i] = -80;
               -79 : lut_out[i] = -80;
               -78 : lut_out[i] = -80;
               -77 : lut_out[i] = -80;
               -76 : lut_out[i] = -80;
               -75 : lut_out[i] = -80;
               -74 : lut_out[i] = -80;
               -73 : lut_out[i] = -64;
               -72 : lut_out[i] = -64;
               -71 : lut_out[i] = -64;
               -70 : lut_out[i] = -64;
               -69 : lut_out[i] = -64;
               -68 : lut_out[i] = -64;
               -67 : lut_out[i] = -64;
               -66 : lut_out[i] = -64;
               -65 : lut_out[i] = -64;
               -64 : lut_out[i] = -64;
               -63 : lut_out[i] = -64;
               -62 : lut_out[i] = -64;
               -61 : lut_out[i] = -64;
               -60 : lut_out[i] = -64;
               -59 : lut_out[i] = -64;
               -58 : lut_out[i] = -64;
               -57 : lut_out[i] = -64;
               -56 : lut_out[i] = -48;
               -55 : lut_out[i] = -48;
               -54 : lut_out[i] = -48;
               -53 : lut_out[i] = -48;
               -52 : lut_out[i] = -48;
               -51 : lut_out[i] = -48;
               -50 : lut_out[i] = -48;
               -49 : lut_out[i] = -48;
               -48 : lut_out[i] = -48;
               -47 : lut_out[i] = -48;
               -46 : lut_out[i] = -48;
               -45 : lut_out[i] = -48;
               -44 : lut_out[i] = -48;
               -43 : lut_out[i] = -48;
               -42 : lut_out[i] = -48;
               -41 : lut_out[i] = -48;
               -40 : lut_out[i] = -32;
               -39 : lut_out[i] = -32;
               -38 : lut_out[i] = -32;
               -37 : lut_out[i] = -32;
               -36 : lut_out[i] = -32;
               -35 : lut_out[i] = -32;
               -34 : lut_out[i] = -32;
               -33 : lut_out[i] = -32;
               -32 : lut_out[i] = -32;
               -31 : lut_out[i] = -32;
               -30 : lut_out[i] = -32;
               -29 : lut_out[i] = -32;
               -28 : lut_out[i] = -32;
               -27 : lut_out[i] = -32;
               -26 : lut_out[i] = -32;
               -25 : lut_out[i] = -32;
               -24 : lut_out[i] = -16;
               -23 : lut_out[i] = -16;
               -22 : lut_out[i] = -16;
               -21 : lut_out[i] = -16;
               -20 : lut_out[i] = -16;
               -19 : lut_out[i] = -16;
               -18 : lut_out[i] = -16;
               -17 : lut_out[i] = -16;
               -16 : lut_out[i] = -16;
               -15 : lut_out[i] = -16;
               -14 : lut_out[i] = -16;
               -13 : lut_out[i] = -16;
               -12 : lut_out[i] = -16;
               -11 : lut_out[i] = -16;
               -10 : lut_out[i] = -16;
               -9 : lut_out[i] = -16;
               -8 : lut_out[i] = 0;
               -7 : lut_out[i] = 0;
               -6 : lut_out[i] = 0;
               -5 : lut_out[i] = 0;
               -4 : lut_out[i] = 0;
               -3 : lut_out[i] = 0;
               -2 : lut_out[i] = 0;
               -1 : lut_out[i] = 0;
               0 : lut_out[i] = 0;
               1 : lut_out[i] = 0;
               2 : lut_out[i] = 0;
               3 : lut_out[i] = 0;
               4 : lut_out[i] = 0;
               5 : lut_out[i] = 0;
               6 : lut_out[i] = 0;
               7 : lut_out[i] = 0;
               8 : lut_out[i] = 0;
               9 : lut_out[i] = 16;
               10 : lut_out[i] = 16;
               11 : lut_out[i] = 16;
               12 : lut_out[i] = 16;
               13 : lut_out[i] = 16;
               14 : lut_out[i] = 16;
               15 : lut_out[i] = 16;
               16 : lut_out[i] = 16;
               17 : lut_out[i] = 16;
               18 : lut_out[i] = 16;
               19 : lut_out[i] = 16;
               20 : lut_out[i] = 16;
               21 : lut_out[i] = 16;
               22 : lut_out[i] = 16;
               23 : lut_out[i] = 16;
               24 : lut_out[i] = 16;
               25 : lut_out[i] = 32;
               26 : lut_out[i] = 32;
               27 : lut_out[i] = 32;
               28 : lut_out[i] = 32;
               29 : lut_out[i] = 32;
               30 : lut_out[i] = 32;
               31 : lut_out[i] = 32;
               32 : lut_out[i] = 32;
               33 : lut_out[i] = 32;
               34 : lut_out[i] = 32;
               35 : lut_out[i] = 32;
               36 : lut_out[i] = 32;
               37 : lut_out[i] = 32;
               38 : lut_out[i] = 32;
               39 : lut_out[i] = 32;
               40 : lut_out[i] = 32;
               41 : lut_out[i] = 48;
               42 : lut_out[i] = 48;
               43 : lut_out[i] = 48;
               44 : lut_out[i] = 48;
               45 : lut_out[i] = 48;
               46 : lut_out[i] = 48;
               47 : lut_out[i] = 48;
               48 : lut_out[i] = 48;
               49 : lut_out[i] = 48;
               50 : lut_out[i] = 48;
               51 : lut_out[i] = 48;
               52 : lut_out[i] = 48;
               53 : lut_out[i] = 48;
               54 : lut_out[i] = 48;
               55 : lut_out[i] = 48;
               56 : lut_out[i] = 48;
               57 : lut_out[i] = 64;
               58 : lut_out[i] = 64;
               59 : lut_out[i] = 64;
               60 : lut_out[i] = 64;
               61 : lut_out[i] = 64;
               62 : lut_out[i] = 64;
               63 : lut_out[i] = 64;
               64 : lut_out[i] = 64;
               65 : lut_out[i] = 64;
               66 : lut_out[i] = 64;
               67 : lut_out[i] = 64;
               68 : lut_out[i] = 64;
               69 : lut_out[i] = 64;
               70 : lut_out[i] = 64;
               71 : lut_out[i] = 64;
               72 : lut_out[i] = 64;
               73 : lut_out[i] = 64;
               74 : lut_out[i] = 80;
               75 : lut_out[i] = 80;
               76 : lut_out[i] = 80;
               77 : lut_out[i] = 80;
               78 : lut_out[i] = 80;
               79 : lut_out[i] = 80;
               80 : lut_out[i] = 80;
               81 : lut_out[i] = 80;
               82 : lut_out[i] = 80;
               83 : lut_out[i] = 80;
               84 : lut_out[i] = 80;
               85 : lut_out[i] = 80;
               86 : lut_out[i] = 80;
               87 : lut_out[i] = 80;
               88 : lut_out[i] = 80;
               89 : lut_out[i] = 80;
               90 : lut_out[i] = 80;
               91 : lut_out[i] = 80;
               92 : lut_out[i] = 96;
               93 : lut_out[i] = 96;
               94 : lut_out[i] = 96;
               95 : lut_out[i] = 96;
               96 : lut_out[i] = 96;
               97 : lut_out[i] = 96;
               98 : lut_out[i] = 96;
               99 : lut_out[i] = 96;
               100 : lut_out[i] = 96;
               101 : lut_out[i] = 96;
               102 : lut_out[i] = 96;
               103 : lut_out[i] = 96;
               104 : lut_out[i] = 96;
               105 : lut_out[i] = 96;
               106 : lut_out[i] = 96;
               107 : lut_out[i] = 96;
               108 : lut_out[i] = 96;
               109 : lut_out[i] = 96;
               110 : lut_out[i] = 96;
               111 : lut_out[i] = 112;
               112 : lut_out[i] = 112;
               113 : lut_out[i] = 112;
               114 : lut_out[i] = 112;
               115 : lut_out[i] = 112;
               116 : lut_out[i] = 112;
               117 : lut_out[i] = 112;
               118 : lut_out[i] = 112;
               119 : lut_out[i] = 112;
               120 : lut_out[i] = 112;
               121 : lut_out[i] = 112;
               122 : lut_out[i] = 112;
               123 : lut_out[i] = 112;
               124 : lut_out[i] = 112;
               125 : lut_out[i] = 112;
               126 : lut_out[i] = 112;
               127 : lut_out[i] = 112;
               128 : lut_out[i] = 112;
               129 : lut_out[i] = 112;
               130 : lut_out[i] = 112;
               131 : lut_out[i] = 128;
               132 : lut_out[i] = 128;
               133 : lut_out[i] = 128;
               134 : lut_out[i] = 128;
               135 : lut_out[i] = 128;
               136 : lut_out[i] = 128;
               137 : lut_out[i] = 128;
               138 : lut_out[i] = 128;
               139 : lut_out[i] = 128;
               140 : lut_out[i] = 128;
               141 : lut_out[i] = 128;
               142 : lut_out[i] = 128;
               143 : lut_out[i] = 128;
               144 : lut_out[i] = 128;
               145 : lut_out[i] = 128;
               146 : lut_out[i] = 128;
               147 : lut_out[i] = 128;
               148 : lut_out[i] = 128;
               149 : lut_out[i] = 128;
               150 : lut_out[i] = 128;
               151 : lut_out[i] = 128;
               152 : lut_out[i] = 144;
               153 : lut_out[i] = 144;
               154 : lut_out[i] = 144;
               155 : lut_out[i] = 144;
               156 : lut_out[i] = 144;
               157 : lut_out[i] = 144;
               158 : lut_out[i] = 144;
               159 : lut_out[i] = 144;
               160 : lut_out[i] = 144;
               161 : lut_out[i] = 144;
               162 : lut_out[i] = 144;
               163 : lut_out[i] = 144;
               164 : lut_out[i] = 144;
               165 : lut_out[i] = 144;
               166 : lut_out[i] = 144;
               167 : lut_out[i] = 144;
               168 : lut_out[i] = 144;
               169 : lut_out[i] = 144;
               170 : lut_out[i] = 144;
               171 : lut_out[i] = 144;
               172 : lut_out[i] = 144;
               173 : lut_out[i] = 144;
               174 : lut_out[i] = 144;
               175 : lut_out[i] = 160;
               176 : lut_out[i] = 160;
               177 : lut_out[i] = 160;
               178 : lut_out[i] = 160;
               179 : lut_out[i] = 160;
               180 : lut_out[i] = 160;
               181 : lut_out[i] = 160;
               182 : lut_out[i] = 160;
               183 : lut_out[i] = 160;
               184 : lut_out[i] = 160;
               185 : lut_out[i] = 160;
               186 : lut_out[i] = 160;
               187 : lut_out[i] = 160;
               188 : lut_out[i] = 160;
               189 : lut_out[i] = 160;
               190 : lut_out[i] = 160;
               191 : lut_out[i] = 160;
               192 : lut_out[i] = 160;
               193 : lut_out[i] = 160;
               194 : lut_out[i] = 160;
               195 : lut_out[i] = 160;
               196 : lut_out[i] = 160;
               197 : lut_out[i] = 160;
               198 : lut_out[i] = 160;
               199 : lut_out[i] = 160;
               200 : lut_out[i] = 160;
               201 : lut_out[i] = 160;
               202 : lut_out[i] = 176;
               203 : lut_out[i] = 176;
               204 : lut_out[i] = 176;
               205 : lut_out[i] = 176;
               206 : lut_out[i] = 176;
               207 : lut_out[i] = 176;
               208 : lut_out[i] = 176;
               209 : lut_out[i] = 176;
               210 : lut_out[i] = 176;
               211 : lut_out[i] = 176;
               212 : lut_out[i] = 176;
               213 : lut_out[i] = 176;
               214 : lut_out[i] = 176;
               215 : lut_out[i] = 176;
               216 : lut_out[i] = 176;
               217 : lut_out[i] = 176;
               218 : lut_out[i] = 176;
               219 : lut_out[i] = 176;
               220 : lut_out[i] = 176;
               221 : lut_out[i] = 176;
               222 : lut_out[i] = 176;
               223 : lut_out[i] = 176;
               224 : lut_out[i] = 176;
               225 : lut_out[i] = 176;
               226 : lut_out[i] = 176;
               227 : lut_out[i] = 176;
               228 : lut_out[i] = 176;
               229 : lut_out[i] = 176;
               230 : lut_out[i] = 176;
               231 : lut_out[i] = 176;
               232 : lut_out[i] = 192;
               233 : lut_out[i] = 192;
               234 : lut_out[i] = 192;
               235 : lut_out[i] = 192;
               236 : lut_out[i] = 192;
               237 : lut_out[i] = 192;
               238 : lut_out[i] = 192;
               239 : lut_out[i] = 192;
               240 : lut_out[i] = 192;
               241 : lut_out[i] = 192;
               242 : lut_out[i] = 192;
               243 : lut_out[i] = 192;
               244 : lut_out[i] = 192;
               245 : lut_out[i] = 192;
               246 : lut_out[i] = 192;
               247 : lut_out[i] = 192;
               248 : lut_out[i] = 192;
               249 : lut_out[i] = 192;
               250 : lut_out[i] = 192;
               251 : lut_out[i] = 192;
               252 : lut_out[i] = 192;
               253 : lut_out[i] = 192;
               254 : lut_out[i] = 192;
               255 : lut_out[i] = 192;
               256 : lut_out[i] = 192;
               257 : lut_out[i] = 192;
               258 : lut_out[i] = 192;
               259 : lut_out[i] = 192;
               260 : lut_out[i] = 192;
               261 : lut_out[i] = 192;
               262 : lut_out[i] = 192;
               263 : lut_out[i] = 192;
               264 : lut_out[i] = 192;
               265 : lut_out[i] = 192;
               266 : lut_out[i] = 192;
               267 : lut_out[i] = 192;
               268 : lut_out[i] = 192;
               269 : lut_out[i] = 208;
               270 : lut_out[i] = 208;
               271 : lut_out[i] = 208;
               272 : lut_out[i] = 208;
               273 : lut_out[i] = 208;
               274 : lut_out[i] = 208;
               275 : lut_out[i] = 208;
               276 : lut_out[i] = 208;
               277 : lut_out[i] = 208;
               278 : lut_out[i] = 208;
               279 : lut_out[i] = 208;
               280 : lut_out[i] = 208;
               281 : lut_out[i] = 208;
               282 : lut_out[i] = 208;
               283 : lut_out[i] = 208;
               284 : lut_out[i] = 208;
               285 : lut_out[i] = 208;
               286 : lut_out[i] = 208;
               287 : lut_out[i] = 208;
               288 : lut_out[i] = 208;
               289 : lut_out[i] = 208;
               290 : lut_out[i] = 208;
               291 : lut_out[i] = 208;
               292 : lut_out[i] = 208;
               293 : lut_out[i] = 208;
               294 : lut_out[i] = 208;
               295 : lut_out[i] = 208;
               296 : lut_out[i] = 208;
               297 : lut_out[i] = 208;
               298 : lut_out[i] = 208;
               299 : lut_out[i] = 208;
               300 : lut_out[i] = 208;
               301 : lut_out[i] = 208;
               302 : lut_out[i] = 208;
               303 : lut_out[i] = 208;
               304 : lut_out[i] = 208;
               305 : lut_out[i] = 208;
               306 : lut_out[i] = 208;
               307 : lut_out[i] = 208;
               308 : lut_out[i] = 208;
               309 : lut_out[i] = 208;
               310 : lut_out[i] = 208;
               311 : lut_out[i] = 208;
               312 : lut_out[i] = 208;
               313 : lut_out[i] = 208;
               314 : lut_out[i] = 208;
               315 : lut_out[i] = 208;
               316 : lut_out[i] = 224;
               317 : lut_out[i] = 224;
               318 : lut_out[i] = 224;
               319 : lut_out[i] = 224;
               320 : lut_out[i] = 224;
               321 : lut_out[i] = 224;
               322 : lut_out[i] = 224;
               323 : lut_out[i] = 224;
               324 : lut_out[i] = 224;
               325 : lut_out[i] = 224;
               326 : lut_out[i] = 224;
               327 : lut_out[i] = 224;
               328 : lut_out[i] = 224;
               329 : lut_out[i] = 224;
               330 : lut_out[i] = 224;
               331 : lut_out[i] = 224;
               332 : lut_out[i] = 224;
               333 : lut_out[i] = 224;
               334 : lut_out[i] = 224;
               335 : lut_out[i] = 224;
               336 : lut_out[i] = 224;
               337 : lut_out[i] = 224;
               338 : lut_out[i] = 224;
               339 : lut_out[i] = 224;
               340 : lut_out[i] = 224;
               341 : lut_out[i] = 224;
               342 : lut_out[i] = 224;
               343 : lut_out[i] = 224;
               344 : lut_out[i] = 224;
               345 : lut_out[i] = 224;
               346 : lut_out[i] = 224;
               347 : lut_out[i] = 224;
               348 : lut_out[i] = 224;
               349 : lut_out[i] = 224;
               350 : lut_out[i] = 224;
               351 : lut_out[i] = 224;
               352 : lut_out[i] = 224;
               353 : lut_out[i] = 224;
               354 : lut_out[i] = 224;
               355 : lut_out[i] = 224;
               356 : lut_out[i] = 224;
               357 : lut_out[i] = 224;
               358 : lut_out[i] = 224;
               359 : lut_out[i] = 224;
               360 : lut_out[i] = 224;
               361 : lut_out[i] = 224;
               362 : lut_out[i] = 224;
               363 : lut_out[i] = 224;
               364 : lut_out[i] = 224;
               365 : lut_out[i] = 224;
               366 : lut_out[i] = 224;
               367 : lut_out[i] = 224;
               368 : lut_out[i] = 224;
               369 : lut_out[i] = 224;
               370 : lut_out[i] = 224;
               371 : lut_out[i] = 224;
               372 : lut_out[i] = 224;
               373 : lut_out[i] = 224;
               374 : lut_out[i] = 224;
               375 : lut_out[i] = 224;
               376 : lut_out[i] = 224;
               377 : lut_out[i] = 224;
               378 : lut_out[i] = 224;
               379 : lut_out[i] = 224;
               380 : lut_out[i] = 224;
               381 : lut_out[i] = 224;
               382 : lut_out[i] = 224;
               383 : lut_out[i] = 224;
               384 : lut_out[i] = 224;
               385 : lut_out[i] = 224;
               386 : lut_out[i] = 240;
               387 : lut_out[i] = 240;
               388 : lut_out[i] = 240;
               389 : lut_out[i] = 240;
               390 : lut_out[i] = 240;
               391 : lut_out[i] = 240;
               392 : lut_out[i] = 240;
               393 : lut_out[i] = 240;
               394 : lut_out[i] = 240;
               395 : lut_out[i] = 240;
               396 : lut_out[i] = 240;
               397 : lut_out[i] = 240;
               398 : lut_out[i] = 240;
               399 : lut_out[i] = 240;
               400 : lut_out[i] = 240;
               401 : lut_out[i] = 240;
               402 : lut_out[i] = 240;
               403 : lut_out[i] = 240;
               404 : lut_out[i] = 240;
               405 : lut_out[i] = 240;
               406 : lut_out[i] = 240;
               407 : lut_out[i] = 240;
               408 : lut_out[i] = 240;
               409 : lut_out[i] = 240;
               410 : lut_out[i] = 240;
               411 : lut_out[i] = 240;
               412 : lut_out[i] = 240;
               413 : lut_out[i] = 240;
               414 : lut_out[i] = 240;
               415 : lut_out[i] = 240;
               416 : lut_out[i] = 240;
               417 : lut_out[i] = 240;
               418 : lut_out[i] = 240;
               419 : lut_out[i] = 240;
               420 : lut_out[i] = 240;
               421 : lut_out[i] = 240;
               422 : lut_out[i] = 240;
               423 : lut_out[i] = 240;
               424 : lut_out[i] = 240;
               425 : lut_out[i] = 240;
               426 : lut_out[i] = 240;
               427 : lut_out[i] = 240;
               428 : lut_out[i] = 240;
               429 : lut_out[i] = 240;
               430 : lut_out[i] = 240;
               431 : lut_out[i] = 240;
               432 : lut_out[i] = 240;
               433 : lut_out[i] = 240;
               434 : lut_out[i] = 240;
               435 : lut_out[i] = 240;
               436 : lut_out[i] = 240;
               437 : lut_out[i] = 240;
               438 : lut_out[i] = 240;
               439 : lut_out[i] = 240;
               440 : lut_out[i] = 240;
               441 : lut_out[i] = 240;
               442 : lut_out[i] = 240;
               443 : lut_out[i] = 240;
               444 : lut_out[i] = 240;
               445 : lut_out[i] = 240;
               446 : lut_out[i] = 240;
               447 : lut_out[i] = 240;
               448 : lut_out[i] = 240;
               449 : lut_out[i] = 240;
               450 : lut_out[i] = 240;
               451 : lut_out[i] = 240;
               452 : lut_out[i] = 240;
               453 : lut_out[i] = 240;
               454 : lut_out[i] = 240;
               455 : lut_out[i] = 240;
               456 : lut_out[i] = 240;
               457 : lut_out[i] = 240;
               458 : lut_out[i] = 240;
               459 : lut_out[i] = 240;
               460 : lut_out[i] = 240;
               461 : lut_out[i] = 240;
               462 : lut_out[i] = 240;
               463 : lut_out[i] = 240;
               464 : lut_out[i] = 240;
               465 : lut_out[i] = 240;
               466 : lut_out[i] = 240;
               467 : lut_out[i] = 240;
               468 : lut_out[i] = 240;
               469 : lut_out[i] = 240;
               470 : lut_out[i] = 240;
               471 : lut_out[i] = 240;
               472 : lut_out[i] = 240;
               473 : lut_out[i] = 240;
               474 : lut_out[i] = 240;
               475 : lut_out[i] = 240;
               476 : lut_out[i] = 240;
               477 : lut_out[i] = 240;
               478 : lut_out[i] = 240;
               479 : lut_out[i] = 240;
               480 : lut_out[i] = 240;
               481 : lut_out[i] = 240;
               482 : lut_out[i] = 240;
               483 : lut_out[i] = 240;
               484 : lut_out[i] = 240;
               485 : lut_out[i] = 240;
               486 : lut_out[i] = 240;
               487 : lut_out[i] = 240;
               488 : lut_out[i] = 240;
               489 : lut_out[i] = 240;
               490 : lut_out[i] = 240;
               491 : lut_out[i] = 240;
               492 : lut_out[i] = 240;
               493 : lut_out[i] = 240;
               494 : lut_out[i] = 240;
               495 : lut_out[i] = 240;
               496 : lut_out[i] = 240;
               497 : lut_out[i] = 240;
               498 : lut_out[i] = 240;
               499 : lut_out[i] = 240;
               500 : lut_out[i] = 240;
               501 : lut_out[i] = 240;
               502 : lut_out[i] = 240;
               503 : lut_out[i] = 240;
               504 : lut_out[i] = 240;
               505 : lut_out[i] = 240;
               506 : lut_out[i] = 240;
               507 : lut_out[i] = 240;
               508 : lut_out[i] = 240;
               509 : lut_out[i] = 240;
               510 : lut_out[i] = 240;
               511 : lut_out[i] = 240;
               512 : lut_out[i] = 240;
               513 : lut_out[i] = 240;
               514 : lut_out[i] = 240;
               515 : lut_out[i] = 240;
               516 : lut_out[i] = 240;
               517 : lut_out[i] = 240;
               518 : lut_out[i] = 240;
               519 : lut_out[i] = 240;
               520 : lut_out[i] = 240;
               521 : lut_out[i] = 240;
               522 : lut_out[i] = 240;
               523 : lut_out[i] = 240;
               524 : lut_out[i] = 240;
               525 : lut_out[i] = 240;
               526 : lut_out[i] = 240;
               527 : lut_out[i] = 240;
               528 : lut_out[i] = 240;
               529 : lut_out[i] = 240;
               530 : lut_out[i] = 240;
               default: lut_out[i] = 0;
            endcase
         end
      end
   end
   
endmodule
