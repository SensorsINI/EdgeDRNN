//-----------------------------------------------------
// Logistic Sigmoid LUT (Q7.8 INPUT & Q0.8 lut_outPUT)
// Design Name : sigmoid_lut.sv
// File Name   : sigmoid_lut.sv
// 
//-----------------------------------------------------
module sigmoid_lut #(
   NUM_PE     = 1,
   ACT_INT_BW = 8,
   ACT_FRA_BW = 8
   )(
   input  logic signed [NUM_PE-1:0][ACT_INT_BW+ACT_FRA_BW-1:0] in,
   output logic signed [NUM_PE-1:0][ACT_INT_BW+ACT_FRA_BW-1:0] out 
   );
   
   localparam ACT_BW = ACT_INT_BW + ACT_FRA_BW;
   logic signed [NUM_PE-1:0][ACT_BW-1:0] lut_in;
   logic signed [NUM_PE-1:0][ACT_BW-1:0] lut_out;
   
   assign out = lut_out;

   always_comb begin
      for (int unsigned i = 0; i < NUM_PE; i = i + 1) begin
         lut_out[i] = '0;
         lut_in[i] = in[i];
         if ($signed(in[i]) > 879) begin // 2047
            lut_out[i] = $signed(256);
         end else if ($signed(in[i]) < -879) begin //-2048
            lut_out[i] = $signed(0);
         end else begin
            case($signed(lut_in[i]))
               -879 : lut_out[i] = 16;
               -878 : lut_out[i] = 16;
               -877 : lut_out[i] = 16;
               -876 : lut_out[i] = 16;
               -875 : lut_out[i] = 16;
               -874 : lut_out[i] = 16;
               -873 : lut_out[i] = 16;
               -872 : lut_out[i] = 16;
               -871 : lut_out[i] = 16;
               -870 : lut_out[i] = 16;
               -869 : lut_out[i] = 16;
               -868 : lut_out[i] = 16;
               -867 : lut_out[i] = 16;
               -866 : lut_out[i] = 16;
               -865 : lut_out[i] = 16;
               -864 : lut_out[i] = 16;
               -863 : lut_out[i] = 16;
               -862 : lut_out[i] = 16;
               -861 : lut_out[i] = 16;
               -860 : lut_out[i] = 16;
               -859 : lut_out[i] = 16;
               -858 : lut_out[i] = 16;
               -857 : lut_out[i] = 16;
               -856 : lut_out[i] = 16;
               -855 : lut_out[i] = 16;
               -854 : lut_out[i] = 16;
               -853 : lut_out[i] = 16;
               -852 : lut_out[i] = 16;
               -851 : lut_out[i] = 16;
               -850 : lut_out[i] = 16;
               -849 : lut_out[i] = 16;
               -848 : lut_out[i] = 16;
               -847 : lut_out[i] = 16;
               -846 : lut_out[i] = 16;
               -845 : lut_out[i] = 16;
               -844 : lut_out[i] = 16;
               -843 : lut_out[i] = 16;
               -842 : lut_out[i] = 16;
               -841 : lut_out[i] = 16;
               -840 : lut_out[i] = 16;
               -839 : lut_out[i] = 16;
               -838 : lut_out[i] = 16;
               -837 : lut_out[i] = 16;
               -836 : lut_out[i] = 16;
               -835 : lut_out[i] = 16;
               -834 : lut_out[i] = 16;
               -833 : lut_out[i] = 16;
               -832 : lut_out[i] = 16;
               -831 : lut_out[i] = 16;
               -830 : lut_out[i] = 16;
               -829 : lut_out[i] = 16;
               -828 : lut_out[i] = 16;
               -827 : lut_out[i] = 16;
               -826 : lut_out[i] = 16;
               -825 : lut_out[i] = 16;
               -824 : lut_out[i] = 16;
               -823 : lut_out[i] = 16;
               -822 : lut_out[i] = 16;
               -821 : lut_out[i] = 16;
               -820 : lut_out[i] = 16;
               -819 : lut_out[i] = 16;
               -818 : lut_out[i] = 16;
               -817 : lut_out[i] = 16;
               -816 : lut_out[i] = 16;
               -815 : lut_out[i] = 16;
               -814 : lut_out[i] = 16;
               -813 : lut_out[i] = 16;
               -812 : lut_out[i] = 16;
               -811 : lut_out[i] = 16;
               -810 : lut_out[i] = 16;
               -809 : lut_out[i] = 16;
               -808 : lut_out[i] = 16;
               -807 : lut_out[i] = 16;
               -806 : lut_out[i] = 16;
               -805 : lut_out[i] = 16;
               -804 : lut_out[i] = 16;
               -803 : lut_out[i] = 16;
               -802 : lut_out[i] = 16;
               -801 : lut_out[i] = 16;
               -800 : lut_out[i] = 16;
               -799 : lut_out[i] = 16;
               -798 : lut_out[i] = 16;
               -797 : lut_out[i] = 16;
               -796 : lut_out[i] = 16;
               -795 : lut_out[i] = 16;
               -794 : lut_out[i] = 16;
               -793 : lut_out[i] = 16;
               -792 : lut_out[i] = 16;
               -791 : lut_out[i] = 16;
               -790 : lut_out[i] = 16;
               -789 : lut_out[i] = 16;
               -788 : lut_out[i] = 16;
               -787 : lut_out[i] = 16;
               -786 : lut_out[i] = 16;
               -785 : lut_out[i] = 16;
               -784 : lut_out[i] = 16;
               -783 : lut_out[i] = 16;
               -782 : lut_out[i] = 16;
               -781 : lut_out[i] = 16;
               -780 : lut_out[i] = 16;
               -779 : lut_out[i] = 16;
               -778 : lut_out[i] = 16;
               -777 : lut_out[i] = 16;
               -776 : lut_out[i] = 16;
               -775 : lut_out[i] = 16;
               -774 : lut_out[i] = 16;
               -773 : lut_out[i] = 16;
               -772 : lut_out[i] = 16;
               -771 : lut_out[i] = 16;
               -770 : lut_out[i] = 16;
               -769 : lut_out[i] = 16;
               -768 : lut_out[i] = 16;
               -767 : lut_out[i] = 16;
               -766 : lut_out[i] = 16;
               -765 : lut_out[i] = 16;
               -764 : lut_out[i] = 16;
               -763 : lut_out[i] = 16;
               -762 : lut_out[i] = 16;
               -761 : lut_out[i] = 16;
               -760 : lut_out[i] = 16;
               -759 : lut_out[i] = 16;
               -758 : lut_out[i] = 16;
               -757 : lut_out[i] = 16;
               -756 : lut_out[i] = 16;
               -755 : lut_out[i] = 16;
               -754 : lut_out[i] = 16;
               -753 : lut_out[i] = 16;
               -752 : lut_out[i] = 16;
               -751 : lut_out[i] = 16;
               -750 : lut_out[i] = 16;
               -749 : lut_out[i] = 16;
               -748 : lut_out[i] = 16;
               -747 : lut_out[i] = 16;
               -746 : lut_out[i] = 16;
               -745 : lut_out[i] = 16;
               -744 : lut_out[i] = 16;
               -743 : lut_out[i] = 16;
               -742 : lut_out[i] = 16;
               -741 : lut_out[i] = 16;
               -740 : lut_out[i] = 16;
               -739 : lut_out[i] = 16;
               -738 : lut_out[i] = 16;
               -737 : lut_out[i] = 16;
               -736 : lut_out[i] = 16;
               -735 : lut_out[i] = 16;
               -734 : lut_out[i] = 16;
               -733 : lut_out[i] = 16;
               -732 : lut_out[i] = 16;
               -731 : lut_out[i] = 16;
               -730 : lut_out[i] = 16;
               -729 : lut_out[i] = 16;
               -728 : lut_out[i] = 16;
               -727 : lut_out[i] = 16;
               -726 : lut_out[i] = 16;
               -725 : lut_out[i] = 16;
               -724 : lut_out[i] = 16;
               -723 : lut_out[i] = 16;
               -722 : lut_out[i] = 16;
               -721 : lut_out[i] = 16;
               -720 : lut_out[i] = 16;
               -719 : lut_out[i] = 16;
               -718 : lut_out[i] = 16;
               -717 : lut_out[i] = 16;
               -716 : lut_out[i] = 16;
               -715 : lut_out[i] = 16;
               -714 : lut_out[i] = 16;
               -713 : lut_out[i] = 16;
               -712 : lut_out[i] = 16;
               -711 : lut_out[i] = 16;
               -710 : lut_out[i] = 16;
               -709 : lut_out[i] = 16;
               -708 : lut_out[i] = 16;
               -707 : lut_out[i] = 16;
               -706 : lut_out[i] = 16;
               -705 : lut_out[i] = 16;
               -704 : lut_out[i] = 16;
               -703 : lut_out[i] = 16;
               -702 : lut_out[i] = 16;
               -701 : lut_out[i] = 16;
               -700 : lut_out[i] = 16;
               -699 : lut_out[i] = 16;
               -698 : lut_out[i] = 16;
               -697 : lut_out[i] = 16;
               -696 : lut_out[i] = 16;
               -695 : lut_out[i] = 16;
               -694 : lut_out[i] = 16;
               -693 : lut_out[i] = 16;
               -692 : lut_out[i] = 16;
               -691 : lut_out[i] = 16;
               -690 : lut_out[i] = 16;
               -689 : lut_out[i] = 16;
               -688 : lut_out[i] = 16;
               -687 : lut_out[i] = 16;
               -686 : lut_out[i] = 16;
               -685 : lut_out[i] = 16;
               -684 : lut_out[i] = 16;
               -683 : lut_out[i] = 16;
               -682 : lut_out[i] = 16;
               -681 : lut_out[i] = 16;
               -680 : lut_out[i] = 16;
               -679 : lut_out[i] = 16;
               -678 : lut_out[i] = 16;
               -677 : lut_out[i] = 16;
               -676 : lut_out[i] = 16;
               -675 : lut_out[i] = 16;
               -674 : lut_out[i] = 16;
               -673 : lut_out[i] = 16;
               -672 : lut_out[i] = 16;
               -671 : lut_out[i] = 16;
               -670 : lut_out[i] = 16;
               -669 : lut_out[i] = 16;
               -668 : lut_out[i] = 16;
               -667 : lut_out[i] = 16;
               -666 : lut_out[i] = 16;
               -665 : lut_out[i] = 16;
               -664 : lut_out[i] = 16;
               -663 : lut_out[i] = 16;
               -662 : lut_out[i] = 16;
               -661 : lut_out[i] = 16;
               -660 : lut_out[i] = 16;
               -659 : lut_out[i] = 16;
               -658 : lut_out[i] = 16;
               -657 : lut_out[i] = 16;
               -656 : lut_out[i] = 16;
               -655 : lut_out[i] = 16;
               -654 : lut_out[i] = 16;
               -653 : lut_out[i] = 16;
               -652 : lut_out[i] = 16;
               -651 : lut_out[i] = 16;
               -650 : lut_out[i] = 16;
               -649 : lut_out[i] = 16;
               -648 : lut_out[i] = 16;
               -647 : lut_out[i] = 16;
               -646 : lut_out[i] = 16;
               -645 : lut_out[i] = 16;
               -644 : lut_out[i] = 16;
               -643 : lut_out[i] = 16;
               -642 : lut_out[i] = 16;
               -641 : lut_out[i] = 16;
               -640 : lut_out[i] = 16;
               -639 : lut_out[i] = 16;
               -638 : lut_out[i] = 16;
               -637 : lut_out[i] = 16;
               -636 : lut_out[i] = 16;
               -635 : lut_out[i] = 16;
               -634 : lut_out[i] = 16;
               -633 : lut_out[i] = 16;
               -632 : lut_out[i] = 16;
               -631 : lut_out[i] = 16;
               -630 : lut_out[i] = 16;
               -629 : lut_out[i] = 16;
               -628 : lut_out[i] = 16;
               -627 : lut_out[i] = 16;
               -626 : lut_out[i] = 16;
               -625 : lut_out[i] = 16;
               -624 : lut_out[i] = 16;
               -623 : lut_out[i] = 16;
               -622 : lut_out[i] = 16;
               -621 : lut_out[i] = 16;
               -620 : lut_out[i] = 16;
               -619 : lut_out[i] = 16;
               -618 : lut_out[i] = 16;
               -617 : lut_out[i] = 16;
               -616 : lut_out[i] = 16;
               -615 : lut_out[i] = 16;
               -614 : lut_out[i] = 16;
               -613 : lut_out[i] = 16;
               -612 : lut_out[i] = 16;
               -611 : lut_out[i] = 16;
               -610 : lut_out[i] = 16;
               -609 : lut_out[i] = 16;
               -608 : lut_out[i] = 16;
               -607 : lut_out[i] = 16;
               -606 : lut_out[i] = 16;
               -605 : lut_out[i] = 16;
               -604 : lut_out[i] = 16;
               -603 : lut_out[i] = 16;
               -602 : lut_out[i] = 16;
               -601 : lut_out[i] = 16;
               -600 : lut_out[i] = 16;
               -599 : lut_out[i] = 16;
               -598 : lut_out[i] = 16;
               -597 : lut_out[i] = 16;
               -596 : lut_out[i] = 16;
               -595 : lut_out[i] = 16;
               -594 : lut_out[i] = 16;
               -593 : lut_out[i] = 16;
               -592 : lut_out[i] = 16;
               -591 : lut_out[i] = 16;
               -590 : lut_out[i] = 16;
               -589 : lut_out[i] = 16;
               -588 : lut_out[i] = 16;
               -587 : lut_out[i] = 16;
               -586 : lut_out[i] = 16;
               -585 : lut_out[i] = 16;
               -584 : lut_out[i] = 16;
               -583 : lut_out[i] = 16;
               -582 : lut_out[i] = 16;
               -581 : lut_out[i] = 16;
               -580 : lut_out[i] = 32;
               -579 : lut_out[i] = 32;
               -578 : lut_out[i] = 32;
               -577 : lut_out[i] = 32;
               -576 : lut_out[i] = 32;
               -575 : lut_out[i] = 32;
               -574 : lut_out[i] = 32;
               -573 : lut_out[i] = 32;
               -572 : lut_out[i] = 32;
               -571 : lut_out[i] = 32;
               -570 : lut_out[i] = 32;
               -569 : lut_out[i] = 32;
               -568 : lut_out[i] = 32;
               -567 : lut_out[i] = 32;
               -566 : lut_out[i] = 32;
               -565 : lut_out[i] = 32;
               -564 : lut_out[i] = 32;
               -563 : lut_out[i] = 32;
               -562 : lut_out[i] = 32;
               -561 : lut_out[i] = 32;
               -560 : lut_out[i] = 32;
               -559 : lut_out[i] = 32;
               -558 : lut_out[i] = 32;
               -557 : lut_out[i] = 32;
               -556 : lut_out[i] = 32;
               -555 : lut_out[i] = 32;
               -554 : lut_out[i] = 32;
               -553 : lut_out[i] = 32;
               -552 : lut_out[i] = 32;
               -551 : lut_out[i] = 32;
               -550 : lut_out[i] = 32;
               -549 : lut_out[i] = 32;
               -548 : lut_out[i] = 32;
               -547 : lut_out[i] = 32;
               -546 : lut_out[i] = 32;
               -545 : lut_out[i] = 32;
               -544 : lut_out[i] = 32;
               -543 : lut_out[i] = 32;
               -542 : lut_out[i] = 32;
               -541 : lut_out[i] = 32;
               -540 : lut_out[i] = 32;
               -539 : lut_out[i] = 32;
               -538 : lut_out[i] = 32;
               -537 : lut_out[i] = 32;
               -536 : lut_out[i] = 32;
               -535 : lut_out[i] = 32;
               -534 : lut_out[i] = 32;
               -533 : lut_out[i] = 32;
               -532 : lut_out[i] = 32;
               -531 : lut_out[i] = 32;
               -530 : lut_out[i] = 32;
               -529 : lut_out[i] = 32;
               -528 : lut_out[i] = 32;
               -527 : lut_out[i] = 32;
               -526 : lut_out[i] = 32;
               -525 : lut_out[i] = 32;
               -524 : lut_out[i] = 32;
               -523 : lut_out[i] = 32;
               -522 : lut_out[i] = 32;
               -521 : lut_out[i] = 32;
               -520 : lut_out[i] = 32;
               -519 : lut_out[i] = 32;
               -518 : lut_out[i] = 32;
               -517 : lut_out[i] = 32;
               -516 : lut_out[i] = 32;
               -515 : lut_out[i] = 32;
               -514 : lut_out[i] = 32;
               -513 : lut_out[i] = 32;
               -512 : lut_out[i] = 32;
               -511 : lut_out[i] = 32;
               -510 : lut_out[i] = 32;
               -509 : lut_out[i] = 32;
               -508 : lut_out[i] = 32;
               -507 : lut_out[i] = 32;
               -506 : lut_out[i] = 32;
               -505 : lut_out[i] = 32;
               -504 : lut_out[i] = 32;
               -503 : lut_out[i] = 32;
               -502 : lut_out[i] = 32;
               -501 : lut_out[i] = 32;
               -500 : lut_out[i] = 32;
               -499 : lut_out[i] = 32;
               -498 : lut_out[i] = 32;
               -497 : lut_out[i] = 32;
               -496 : lut_out[i] = 32;
               -495 : lut_out[i] = 32;
               -494 : lut_out[i] = 32;
               -493 : lut_out[i] = 32;
               -492 : lut_out[i] = 32;
               -491 : lut_out[i] = 32;
               -490 : lut_out[i] = 32;
               -489 : lut_out[i] = 32;
               -488 : lut_out[i] = 32;
               -487 : lut_out[i] = 32;
               -486 : lut_out[i] = 32;
               -485 : lut_out[i] = 32;
               -484 : lut_out[i] = 32;
               -483 : lut_out[i] = 32;
               -482 : lut_out[i] = 32;
               -481 : lut_out[i] = 32;
               -480 : lut_out[i] = 32;
               -479 : lut_out[i] = 32;
               -478 : lut_out[i] = 32;
               -477 : lut_out[i] = 32;
               -476 : lut_out[i] = 32;
               -475 : lut_out[i] = 32;
               -474 : lut_out[i] = 32;
               -473 : lut_out[i] = 32;
               -472 : lut_out[i] = 32;
               -471 : lut_out[i] = 32;
               -470 : lut_out[i] = 32;
               -469 : lut_out[i] = 32;
               -468 : lut_out[i] = 32;
               -467 : lut_out[i] = 32;
               -466 : lut_out[i] = 32;
               -465 : lut_out[i] = 32;
               -464 : lut_out[i] = 32;
               -463 : lut_out[i] = 32;
               -462 : lut_out[i] = 32;
               -461 : lut_out[i] = 32;
               -460 : lut_out[i] = 32;
               -459 : lut_out[i] = 32;
               -458 : lut_out[i] = 32;
               -457 : lut_out[i] = 32;
               -456 : lut_out[i] = 32;
               -455 : lut_out[i] = 32;
               -454 : lut_out[i] = 32;
               -453 : lut_out[i] = 32;
               -452 : lut_out[i] = 32;
               -451 : lut_out[i] = 32;
               -450 : lut_out[i] = 32;
               -449 : lut_out[i] = 32;
               -448 : lut_out[i] = 32;
               -447 : lut_out[i] = 32;
               -446 : lut_out[i] = 32;
               -445 : lut_out[i] = 32;
               -444 : lut_out[i] = 32;
               -443 : lut_out[i] = 32;
               -442 : lut_out[i] = 32;
               -441 : lut_out[i] = 32;
               -440 : lut_out[i] = 32;
               -439 : lut_out[i] = 32;
               -438 : lut_out[i] = 32;
               -437 : lut_out[i] = 32;
               -436 : lut_out[i] = 32;
               -435 : lut_out[i] = 32;
               -434 : lut_out[i] = 32;
               -433 : lut_out[i] = 32;
               -432 : lut_out[i] = 32;
               -431 : lut_out[i] = 48;
               -430 : lut_out[i] = 48;
               -429 : lut_out[i] = 48;
               -428 : lut_out[i] = 48;
               -427 : lut_out[i] = 48;
               -426 : lut_out[i] = 48;
               -425 : lut_out[i] = 48;
               -424 : lut_out[i] = 48;
               -423 : lut_out[i] = 48;
               -422 : lut_out[i] = 48;
               -421 : lut_out[i] = 48;
               -420 : lut_out[i] = 48;
               -419 : lut_out[i] = 48;
               -418 : lut_out[i] = 48;
               -417 : lut_out[i] = 48;
               -416 : lut_out[i] = 48;
               -415 : lut_out[i] = 48;
               -414 : lut_out[i] = 48;
               -413 : lut_out[i] = 48;
               -412 : lut_out[i] = 48;
               -411 : lut_out[i] = 48;
               -410 : lut_out[i] = 48;
               -409 : lut_out[i] = 48;
               -408 : lut_out[i] = 48;
               -407 : lut_out[i] = 48;
               -406 : lut_out[i] = 48;
               -405 : lut_out[i] = 48;
               -404 : lut_out[i] = 48;
               -403 : lut_out[i] = 48;
               -402 : lut_out[i] = 48;
               -401 : lut_out[i] = 48;
               -400 : lut_out[i] = 48;
               -399 : lut_out[i] = 48;
               -398 : lut_out[i] = 48;
               -397 : lut_out[i] = 48;
               -396 : lut_out[i] = 48;
               -395 : lut_out[i] = 48;
               -394 : lut_out[i] = 48;
               -393 : lut_out[i] = 48;
               -392 : lut_out[i] = 48;
               -391 : lut_out[i] = 48;
               -390 : lut_out[i] = 48;
               -389 : lut_out[i] = 48;
               -388 : lut_out[i] = 48;
               -387 : lut_out[i] = 48;
               -386 : lut_out[i] = 48;
               -385 : lut_out[i] = 48;
               -384 : lut_out[i] = 48;
               -383 : lut_out[i] = 48;
               -382 : lut_out[i] = 48;
               -381 : lut_out[i] = 48;
               -380 : lut_out[i] = 48;
               -379 : lut_out[i] = 48;
               -378 : lut_out[i] = 48;
               -377 : lut_out[i] = 48;
               -376 : lut_out[i] = 48;
               -375 : lut_out[i] = 48;
               -374 : lut_out[i] = 48;
               -373 : lut_out[i] = 48;
               -372 : lut_out[i] = 48;
               -371 : lut_out[i] = 48;
               -370 : lut_out[i] = 48;
               -369 : lut_out[i] = 48;
               -368 : lut_out[i] = 48;
               -367 : lut_out[i] = 48;
               -366 : lut_out[i] = 48;
               -365 : lut_out[i] = 48;
               -364 : lut_out[i] = 48;
               -363 : lut_out[i] = 48;
               -362 : lut_out[i] = 48;
               -361 : lut_out[i] = 48;
               -360 : lut_out[i] = 48;
               -359 : lut_out[i] = 48;
               -358 : lut_out[i] = 48;
               -357 : lut_out[i] = 48;
               -356 : lut_out[i] = 48;
               -355 : lut_out[i] = 48;
               -354 : lut_out[i] = 48;
               -353 : lut_out[i] = 48;
               -352 : lut_out[i] = 48;
               -351 : lut_out[i] = 48;
               -350 : lut_out[i] = 48;
               -349 : lut_out[i] = 48;
               -348 : lut_out[i] = 48;
               -347 : lut_out[i] = 48;
               -346 : lut_out[i] = 48;
               -345 : lut_out[i] = 48;
               -344 : lut_out[i] = 48;
               -343 : lut_out[i] = 48;
               -342 : lut_out[i] = 48;
               -341 : lut_out[i] = 48;
               -340 : lut_out[i] = 48;
               -339 : lut_out[i] = 48;
               -338 : lut_out[i] = 48;
               -337 : lut_out[i] = 48;
               -336 : lut_out[i] = 48;
               -335 : lut_out[i] = 48;
               -334 : lut_out[i] = 48;
               -333 : lut_out[i] = 48;
               -332 : lut_out[i] = 48;
               -331 : lut_out[i] = 48;
               -330 : lut_out[i] = 48;
               -329 : lut_out[i] = 48;
               -328 : lut_out[i] = 48;
               -327 : lut_out[i] = 48;
               -326 : lut_out[i] = 48;
               -325 : lut_out[i] = 64;
               -324 : lut_out[i] = 64;
               -323 : lut_out[i] = 64;
               -322 : lut_out[i] = 64;
               -321 : lut_out[i] = 64;
               -320 : lut_out[i] = 64;
               -319 : lut_out[i] = 64;
               -318 : lut_out[i] = 64;
               -317 : lut_out[i] = 64;
               -316 : lut_out[i] = 64;
               -315 : lut_out[i] = 64;
               -314 : lut_out[i] = 64;
               -313 : lut_out[i] = 64;
               -312 : lut_out[i] = 64;
               -311 : lut_out[i] = 64;
               -310 : lut_out[i] = 64;
               -309 : lut_out[i] = 64;
               -308 : lut_out[i] = 64;
               -307 : lut_out[i] = 64;
               -306 : lut_out[i] = 64;
               -305 : lut_out[i] = 64;
               -304 : lut_out[i] = 64;
               -303 : lut_out[i] = 64;
               -302 : lut_out[i] = 64;
               -301 : lut_out[i] = 64;
               -300 : lut_out[i] = 64;
               -299 : lut_out[i] = 64;
               -298 : lut_out[i] = 64;
               -297 : lut_out[i] = 64;
               -296 : lut_out[i] = 64;
               -295 : lut_out[i] = 64;
               -294 : lut_out[i] = 64;
               -293 : lut_out[i] = 64;
               -292 : lut_out[i] = 64;
               -291 : lut_out[i] = 64;
               -290 : lut_out[i] = 64;
               -289 : lut_out[i] = 64;
               -288 : lut_out[i] = 64;
               -287 : lut_out[i] = 64;
               -286 : lut_out[i] = 64;
               -285 : lut_out[i] = 64;
               -284 : lut_out[i] = 64;
               -283 : lut_out[i] = 64;
               -282 : lut_out[i] = 64;
               -281 : lut_out[i] = 64;
               -280 : lut_out[i] = 64;
               -279 : lut_out[i] = 64;
               -278 : lut_out[i] = 64;
               -277 : lut_out[i] = 64;
               -276 : lut_out[i] = 64;
               -275 : lut_out[i] = 64;
               -274 : lut_out[i] = 64;
               -273 : lut_out[i] = 64;
               -272 : lut_out[i] = 64;
               -271 : lut_out[i] = 64;
               -270 : lut_out[i] = 64;
               -269 : lut_out[i] = 64;
               -268 : lut_out[i] = 64;
               -267 : lut_out[i] = 64;
               -266 : lut_out[i] = 64;
               -265 : lut_out[i] = 64;
               -264 : lut_out[i] = 64;
               -263 : lut_out[i] = 64;
               -262 : lut_out[i] = 64;
               -261 : lut_out[i] = 64;
               -260 : lut_out[i] = 64;
               -259 : lut_out[i] = 64;
               -258 : lut_out[i] = 64;
               -257 : lut_out[i] = 64;
               -256 : lut_out[i] = 64;
               -255 : lut_out[i] = 64;
               -254 : lut_out[i] = 64;
               -253 : lut_out[i] = 64;
               -252 : lut_out[i] = 64;
               -251 : lut_out[i] = 64;
               -250 : lut_out[i] = 64;
               -249 : lut_out[i] = 64;
               -248 : lut_out[i] = 64;
               -247 : lut_out[i] = 64;
               -246 : lut_out[i] = 64;
               -245 : lut_out[i] = 64;
               -244 : lut_out[i] = 64;
               -243 : lut_out[i] = 64;
               -242 : lut_out[i] = 64;
               -241 : lut_out[i] = 64;
               -240 : lut_out[i] = 80;
               -239 : lut_out[i] = 80;
               -238 : lut_out[i] = 80;
               -237 : lut_out[i] = 80;
               -236 : lut_out[i] = 80;
               -235 : lut_out[i] = 80;
               -234 : lut_out[i] = 80;
               -233 : lut_out[i] = 80;
               -232 : lut_out[i] = 80;
               -231 : lut_out[i] = 80;
               -230 : lut_out[i] = 80;
               -229 : lut_out[i] = 80;
               -228 : lut_out[i] = 80;
               -227 : lut_out[i] = 80;
               -226 : lut_out[i] = 80;
               -225 : lut_out[i] = 80;
               -224 : lut_out[i] = 80;
               -223 : lut_out[i] = 80;
               -222 : lut_out[i] = 80;
               -221 : lut_out[i] = 80;
               -220 : lut_out[i] = 80;
               -219 : lut_out[i] = 80;
               -218 : lut_out[i] = 80;
               -217 : lut_out[i] = 80;
               -216 : lut_out[i] = 80;
               -215 : lut_out[i] = 80;
               -214 : lut_out[i] = 80;
               -213 : lut_out[i] = 80;
               -212 : lut_out[i] = 80;
               -211 : lut_out[i] = 80;
               -210 : lut_out[i] = 80;
               -209 : lut_out[i] = 80;
               -208 : lut_out[i] = 80;
               -207 : lut_out[i] = 80;
               -206 : lut_out[i] = 80;
               -205 : lut_out[i] = 80;
               -204 : lut_out[i] = 80;
               -203 : lut_out[i] = 80;
               -202 : lut_out[i] = 80;
               -201 : lut_out[i] = 80;
               -200 : lut_out[i] = 80;
               -199 : lut_out[i] = 80;
               -198 : lut_out[i] = 80;
               -197 : lut_out[i] = 80;
               -196 : lut_out[i] = 80;
               -195 : lut_out[i] = 80;
               -194 : lut_out[i] = 80;
               -193 : lut_out[i] = 80;
               -192 : lut_out[i] = 80;
               -191 : lut_out[i] = 80;
               -190 : lut_out[i] = 80;
               -189 : lut_out[i] = 80;
               -188 : lut_out[i] = 80;
               -187 : lut_out[i] = 80;
               -186 : lut_out[i] = 80;
               -185 : lut_out[i] = 80;
               -184 : lut_out[i] = 80;
               -183 : lut_out[i] = 80;
               -182 : lut_out[i] = 80;
               -181 : lut_out[i] = 80;
               -180 : lut_out[i] = 80;
               -179 : lut_out[i] = 80;
               -178 : lut_out[i] = 80;
               -177 : lut_out[i] = 80;
               -176 : lut_out[i] = 80;
               -175 : lut_out[i] = 80;
               -174 : lut_out[i] = 80;
               -173 : lut_out[i] = 80;
               -172 : lut_out[i] = 80;
               -171 : lut_out[i] = 80;
               -170 : lut_out[i] = 80;
               -169 : lut_out[i] = 80;
               -168 : lut_out[i] = 80;
               -167 : lut_out[i] = 80;
               -166 : lut_out[i] = 80;
               -165 : lut_out[i] = 96;
               -164 : lut_out[i] = 96;
               -163 : lut_out[i] = 96;
               -162 : lut_out[i] = 96;
               -161 : lut_out[i] = 96;
               -160 : lut_out[i] = 96;
               -159 : lut_out[i] = 96;
               -158 : lut_out[i] = 96;
               -157 : lut_out[i] = 96;
               -156 : lut_out[i] = 96;
               -155 : lut_out[i] = 96;
               -154 : lut_out[i] = 96;
               -153 : lut_out[i] = 96;
               -152 : lut_out[i] = 96;
               -151 : lut_out[i] = 96;
               -150 : lut_out[i] = 96;
               -149 : lut_out[i] = 96;
               -148 : lut_out[i] = 96;
               -147 : lut_out[i] = 96;
               -146 : lut_out[i] = 96;
               -145 : lut_out[i] = 96;
               -144 : lut_out[i] = 96;
               -143 : lut_out[i] = 96;
               -142 : lut_out[i] = 96;
               -141 : lut_out[i] = 96;
               -140 : lut_out[i] = 96;
               -139 : lut_out[i] = 96;
               -138 : lut_out[i] = 96;
               -137 : lut_out[i] = 96;
               -136 : lut_out[i] = 96;
               -135 : lut_out[i] = 96;
               -134 : lut_out[i] = 96;
               -133 : lut_out[i] = 96;
               -132 : lut_out[i] = 96;
               -131 : lut_out[i] = 96;
               -130 : lut_out[i] = 96;
               -129 : lut_out[i] = 96;
               -128 : lut_out[i] = 96;
               -127 : lut_out[i] = 96;
               -126 : lut_out[i] = 96;
               -125 : lut_out[i] = 96;
               -124 : lut_out[i] = 96;
               -123 : lut_out[i] = 96;
               -122 : lut_out[i] = 96;
               -121 : lut_out[i] = 96;
               -120 : lut_out[i] = 96;
               -119 : lut_out[i] = 96;
               -118 : lut_out[i] = 96;
               -117 : lut_out[i] = 96;
               -116 : lut_out[i] = 96;
               -115 : lut_out[i] = 96;
               -114 : lut_out[i] = 96;
               -113 : lut_out[i] = 96;
               -112 : lut_out[i] = 96;
               -111 : lut_out[i] = 96;
               -110 : lut_out[i] = 96;
               -109 : lut_out[i] = 96;
               -108 : lut_out[i] = 96;
               -107 : lut_out[i] = 96;
               -106 : lut_out[i] = 96;
               -105 : lut_out[i] = 96;
               -104 : lut_out[i] = 96;
               -103 : lut_out[i] = 96;
               -102 : lut_out[i] = 96;
               -101 : lut_out[i] = 96;
               -100 : lut_out[i] = 96;
               -99 : lut_out[i] = 96;
               -98 : lut_out[i] = 96;
               -97 : lut_out[i] = 112;
               -96 : lut_out[i] = 112;
               -95 : lut_out[i] = 112;
               -94 : lut_out[i] = 112;
               -93 : lut_out[i] = 112;
               -92 : lut_out[i] = 112;
               -91 : lut_out[i] = 112;
               -90 : lut_out[i] = 112;
               -89 : lut_out[i] = 112;
               -88 : lut_out[i] = 112;
               -87 : lut_out[i] = 112;
               -86 : lut_out[i] = 112;
               -85 : lut_out[i] = 112;
               -84 : lut_out[i] = 112;
               -83 : lut_out[i] = 112;
               -82 : lut_out[i] = 112;
               -81 : lut_out[i] = 112;
               -80 : lut_out[i] = 112;
               -79 : lut_out[i] = 112;
               -78 : lut_out[i] = 112;
               -77 : lut_out[i] = 112;
               -76 : lut_out[i] = 112;
               -75 : lut_out[i] = 112;
               -74 : lut_out[i] = 112;
               -73 : lut_out[i] = 112;
               -72 : lut_out[i] = 112;
               -71 : lut_out[i] = 112;
               -70 : lut_out[i] = 112;
               -69 : lut_out[i] = 112;
               -68 : lut_out[i] = 112;
               -67 : lut_out[i] = 112;
               -66 : lut_out[i] = 112;
               -65 : lut_out[i] = 112;
               -64 : lut_out[i] = 112;
               -63 : lut_out[i] = 112;
               -62 : lut_out[i] = 112;
               -61 : lut_out[i] = 112;
               -60 : lut_out[i] = 112;
               -59 : lut_out[i] = 112;
               -58 : lut_out[i] = 112;
               -57 : lut_out[i] = 112;
               -56 : lut_out[i] = 112;
               -55 : lut_out[i] = 112;
               -54 : lut_out[i] = 112;
               -53 : lut_out[i] = 112;
               -52 : lut_out[i] = 112;
               -51 : lut_out[i] = 112;
               -50 : lut_out[i] = 112;
               -49 : lut_out[i] = 112;
               -48 : lut_out[i] = 112;
               -47 : lut_out[i] = 112;
               -46 : lut_out[i] = 112;
               -45 : lut_out[i] = 112;
               -44 : lut_out[i] = 112;
               -43 : lut_out[i] = 112;
               -42 : lut_out[i] = 112;
               -41 : lut_out[i] = 112;
               -40 : lut_out[i] = 112;
               -39 : lut_out[i] = 112;
               -38 : lut_out[i] = 112;
               -37 : lut_out[i] = 112;
               -36 : lut_out[i] = 112;
               -35 : lut_out[i] = 112;
               -34 : lut_out[i] = 112;
               -33 : lut_out[i] = 112;
               -32 : lut_out[i] = 128;
               -31 : lut_out[i] = 128;
               -30 : lut_out[i] = 128;
               -29 : lut_out[i] = 128;
               -28 : lut_out[i] = 128;
               -27 : lut_out[i] = 128;
               -26 : lut_out[i] = 128;
               -25 : lut_out[i] = 128;
               -24 : lut_out[i] = 128;
               -23 : lut_out[i] = 128;
               -22 : lut_out[i] = 128;
               -21 : lut_out[i] = 128;
               -20 : lut_out[i] = 128;
               -19 : lut_out[i] = 128;
               -18 : lut_out[i] = 128;
               -17 : lut_out[i] = 128;
               -16 : lut_out[i] = 128;
               -15 : lut_out[i] = 128;
               -14 : lut_out[i] = 128;
               -13 : lut_out[i] = 128;
               -12 : lut_out[i] = 128;
               -11 : lut_out[i] = 128;
               -10 : lut_out[i] = 128;
               -9 : lut_out[i] = 128;
               -8 : lut_out[i] = 128;
               -7 : lut_out[i] = 128;
               -6 : lut_out[i] = 128;
               -5 : lut_out[i] = 128;
               -4 : lut_out[i] = 128;
               -3 : lut_out[i] = 128;
               -2 : lut_out[i] = 128;
               -1 : lut_out[i] = 128;
               0 : lut_out[i] = 128;
               1 : lut_out[i] = 128;
               2 : lut_out[i] = 128;
               3 : lut_out[i] = 128;
               4 : lut_out[i] = 128;
               5 : lut_out[i] = 128;
               6 : lut_out[i] = 128;
               7 : lut_out[i] = 128;
               8 : lut_out[i] = 128;
               9 : lut_out[i] = 128;
               10 : lut_out[i] = 128;
               11 : lut_out[i] = 128;
               12 : lut_out[i] = 128;
               13 : lut_out[i] = 128;
               14 : lut_out[i] = 128;
               15 : lut_out[i] = 128;
               16 : lut_out[i] = 128;
               17 : lut_out[i] = 128;
               18 : lut_out[i] = 128;
               19 : lut_out[i] = 128;
               20 : lut_out[i] = 128;
               21 : lut_out[i] = 128;
               22 : lut_out[i] = 128;
               23 : lut_out[i] = 128;
               24 : lut_out[i] = 128;
               25 : lut_out[i] = 128;
               26 : lut_out[i] = 128;
               27 : lut_out[i] = 128;
               28 : lut_out[i] = 128;
               29 : lut_out[i] = 128;
               30 : lut_out[i] = 128;
               31 : lut_out[i] = 128;
               32 : lut_out[i] = 128;
               33 : lut_out[i] = 144;
               34 : lut_out[i] = 144;
               35 : lut_out[i] = 144;
               36 : lut_out[i] = 144;
               37 : lut_out[i] = 144;
               38 : lut_out[i] = 144;
               39 : lut_out[i] = 144;
               40 : lut_out[i] = 144;
               41 : lut_out[i] = 144;
               42 : lut_out[i] = 144;
               43 : lut_out[i] = 144;
               44 : lut_out[i] = 144;
               45 : lut_out[i] = 144;
               46 : lut_out[i] = 144;
               47 : lut_out[i] = 144;
               48 : lut_out[i] = 144;
               49 : lut_out[i] = 144;
               50 : lut_out[i] = 144;
               51 : lut_out[i] = 144;
               52 : lut_out[i] = 144;
               53 : lut_out[i] = 144;
               54 : lut_out[i] = 144;
               55 : lut_out[i] = 144;
               56 : lut_out[i] = 144;
               57 : lut_out[i] = 144;
               58 : lut_out[i] = 144;
               59 : lut_out[i] = 144;
               60 : lut_out[i] = 144;
               61 : lut_out[i] = 144;
               62 : lut_out[i] = 144;
               63 : lut_out[i] = 144;
               64 : lut_out[i] = 144;
               65 : lut_out[i] = 144;
               66 : lut_out[i] = 144;
               67 : lut_out[i] = 144;
               68 : lut_out[i] = 144;
               69 : lut_out[i] = 144;
               70 : lut_out[i] = 144;
               71 : lut_out[i] = 144;
               72 : lut_out[i] = 144;
               73 : lut_out[i] = 144;
               74 : lut_out[i] = 144;
               75 : lut_out[i] = 144;
               76 : lut_out[i] = 144;
               77 : lut_out[i] = 144;
               78 : lut_out[i] = 144;
               79 : lut_out[i] = 144;
               80 : lut_out[i] = 144;
               81 : lut_out[i] = 144;
               82 : lut_out[i] = 144;
               83 : lut_out[i] = 144;
               84 : lut_out[i] = 144;
               85 : lut_out[i] = 144;
               86 : lut_out[i] = 144;
               87 : lut_out[i] = 144;
               88 : lut_out[i] = 144;
               89 : lut_out[i] = 144;
               90 : lut_out[i] = 144;
               91 : lut_out[i] = 144;
               92 : lut_out[i] = 144;
               93 : lut_out[i] = 144;
               94 : lut_out[i] = 144;
               95 : lut_out[i] = 144;
               96 : lut_out[i] = 144;
               97 : lut_out[i] = 144;
               98 : lut_out[i] = 160;
               99 : lut_out[i] = 160;
               100 : lut_out[i] = 160;
               101 : lut_out[i] = 160;
               102 : lut_out[i] = 160;
               103 : lut_out[i] = 160;
               104 : lut_out[i] = 160;
               105 : lut_out[i] = 160;
               106 : lut_out[i] = 160;
               107 : lut_out[i] = 160;
               108 : lut_out[i] = 160;
               109 : lut_out[i] = 160;
               110 : lut_out[i] = 160;
               111 : lut_out[i] = 160;
               112 : lut_out[i] = 160;
               113 : lut_out[i] = 160;
               114 : lut_out[i] = 160;
               115 : lut_out[i] = 160;
               116 : lut_out[i] = 160;
               117 : lut_out[i] = 160;
               118 : lut_out[i] = 160;
               119 : lut_out[i] = 160;
               120 : lut_out[i] = 160;
               121 : lut_out[i] = 160;
               122 : lut_out[i] = 160;
               123 : lut_out[i] = 160;
               124 : lut_out[i] = 160;
               125 : lut_out[i] = 160;
               126 : lut_out[i] = 160;
               127 : lut_out[i] = 160;
               128 : lut_out[i] = 160;
               129 : lut_out[i] = 160;
               130 : lut_out[i] = 160;
               131 : lut_out[i] = 160;
               132 : lut_out[i] = 160;
               133 : lut_out[i] = 160;
               134 : lut_out[i] = 160;
               135 : lut_out[i] = 160;
               136 : lut_out[i] = 160;
               137 : lut_out[i] = 160;
               138 : lut_out[i] = 160;
               139 : lut_out[i] = 160;
               140 : lut_out[i] = 160;
               141 : lut_out[i] = 160;
               142 : lut_out[i] = 160;
               143 : lut_out[i] = 160;
               144 : lut_out[i] = 160;
               145 : lut_out[i] = 160;
               146 : lut_out[i] = 160;
               147 : lut_out[i] = 160;
               148 : lut_out[i] = 160;
               149 : lut_out[i] = 160;
               150 : lut_out[i] = 160;
               151 : lut_out[i] = 160;
               152 : lut_out[i] = 160;
               153 : lut_out[i] = 160;
               154 : lut_out[i] = 160;
               155 : lut_out[i] = 160;
               156 : lut_out[i] = 160;
               157 : lut_out[i] = 160;
               158 : lut_out[i] = 160;
               159 : lut_out[i] = 160;
               160 : lut_out[i] = 160;
               161 : lut_out[i] = 160;
               162 : lut_out[i] = 160;
               163 : lut_out[i] = 160;
               164 : lut_out[i] = 160;
               165 : lut_out[i] = 160;
               166 : lut_out[i] = 176;
               167 : lut_out[i] = 176;
               168 : lut_out[i] = 176;
               169 : lut_out[i] = 176;
               170 : lut_out[i] = 176;
               171 : lut_out[i] = 176;
               172 : lut_out[i] = 176;
               173 : lut_out[i] = 176;
               174 : lut_out[i] = 176;
               175 : lut_out[i] = 176;
               176 : lut_out[i] = 176;
               177 : lut_out[i] = 176;
               178 : lut_out[i] = 176;
               179 : lut_out[i] = 176;
               180 : lut_out[i] = 176;
               181 : lut_out[i] = 176;
               182 : lut_out[i] = 176;
               183 : lut_out[i] = 176;
               184 : lut_out[i] = 176;
               185 : lut_out[i] = 176;
               186 : lut_out[i] = 176;
               187 : lut_out[i] = 176;
               188 : lut_out[i] = 176;
               189 : lut_out[i] = 176;
               190 : lut_out[i] = 176;
               191 : lut_out[i] = 176;
               192 : lut_out[i] = 176;
               193 : lut_out[i] = 176;
               194 : lut_out[i] = 176;
               195 : lut_out[i] = 176;
               196 : lut_out[i] = 176;
               197 : lut_out[i] = 176;
               198 : lut_out[i] = 176;
               199 : lut_out[i] = 176;
               200 : lut_out[i] = 176;
               201 : lut_out[i] = 176;
               202 : lut_out[i] = 176;
               203 : lut_out[i] = 176;
               204 : lut_out[i] = 176;
               205 : lut_out[i] = 176;
               206 : lut_out[i] = 176;
               207 : lut_out[i] = 176;
               208 : lut_out[i] = 176;
               209 : lut_out[i] = 176;
               210 : lut_out[i] = 176;
               211 : lut_out[i] = 176;
               212 : lut_out[i] = 176;
               213 : lut_out[i] = 176;
               214 : lut_out[i] = 176;
               215 : lut_out[i] = 176;
               216 : lut_out[i] = 176;
               217 : lut_out[i] = 176;
               218 : lut_out[i] = 176;
               219 : lut_out[i] = 176;
               220 : lut_out[i] = 176;
               221 : lut_out[i] = 176;
               222 : lut_out[i] = 176;
               223 : lut_out[i] = 176;
               224 : lut_out[i] = 176;
               225 : lut_out[i] = 176;
               226 : lut_out[i] = 176;
               227 : lut_out[i] = 176;
               228 : lut_out[i] = 176;
               229 : lut_out[i] = 176;
               230 : lut_out[i] = 176;
               231 : lut_out[i] = 176;
               232 : lut_out[i] = 176;
               233 : lut_out[i] = 176;
               234 : lut_out[i] = 176;
               235 : lut_out[i] = 176;
               236 : lut_out[i] = 176;
               237 : lut_out[i] = 176;
               238 : lut_out[i] = 176;
               239 : lut_out[i] = 176;
               240 : lut_out[i] = 176;
               241 : lut_out[i] = 192;
               242 : lut_out[i] = 192;
               243 : lut_out[i] = 192;
               244 : lut_out[i] = 192;
               245 : lut_out[i] = 192;
               246 : lut_out[i] = 192;
               247 : lut_out[i] = 192;
               248 : lut_out[i] = 192;
               249 : lut_out[i] = 192;
               250 : lut_out[i] = 192;
               251 : lut_out[i] = 192;
               252 : lut_out[i] = 192;
               253 : lut_out[i] = 192;
               254 : lut_out[i] = 192;
               255 : lut_out[i] = 192;
               256 : lut_out[i] = 192;
               257 : lut_out[i] = 192;
               258 : lut_out[i] = 192;
               259 : lut_out[i] = 192;
               260 : lut_out[i] = 192;
               261 : lut_out[i] = 192;
               262 : lut_out[i] = 192;
               263 : lut_out[i] = 192;
               264 : lut_out[i] = 192;
               265 : lut_out[i] = 192;
               266 : lut_out[i] = 192;
               267 : lut_out[i] = 192;
               268 : lut_out[i] = 192;
               269 : lut_out[i] = 192;
               270 : lut_out[i] = 192;
               271 : lut_out[i] = 192;
               272 : lut_out[i] = 192;
               273 : lut_out[i] = 192;
               274 : lut_out[i] = 192;
               275 : lut_out[i] = 192;
               276 : lut_out[i] = 192;
               277 : lut_out[i] = 192;
               278 : lut_out[i] = 192;
               279 : lut_out[i] = 192;
               280 : lut_out[i] = 192;
               281 : lut_out[i] = 192;
               282 : lut_out[i] = 192;
               283 : lut_out[i] = 192;
               284 : lut_out[i] = 192;
               285 : lut_out[i] = 192;
               286 : lut_out[i] = 192;
               287 : lut_out[i] = 192;
               288 : lut_out[i] = 192;
               289 : lut_out[i] = 192;
               290 : lut_out[i] = 192;
               291 : lut_out[i] = 192;
               292 : lut_out[i] = 192;
               293 : lut_out[i] = 192;
               294 : lut_out[i] = 192;
               295 : lut_out[i] = 192;
               296 : lut_out[i] = 192;
               297 : lut_out[i] = 192;
               298 : lut_out[i] = 192;
               299 : lut_out[i] = 192;
               300 : lut_out[i] = 192;
               301 : lut_out[i] = 192;
               302 : lut_out[i] = 192;
               303 : lut_out[i] = 192;
               304 : lut_out[i] = 192;
               305 : lut_out[i] = 192;
               306 : lut_out[i] = 192;
               307 : lut_out[i] = 192;
               308 : lut_out[i] = 192;
               309 : lut_out[i] = 192;
               310 : lut_out[i] = 192;
               311 : lut_out[i] = 192;
               312 : lut_out[i] = 192;
               313 : lut_out[i] = 192;
               314 : lut_out[i] = 192;
               315 : lut_out[i] = 192;
               316 : lut_out[i] = 192;
               317 : lut_out[i] = 192;
               318 : lut_out[i] = 192;
               319 : lut_out[i] = 192;
               320 : lut_out[i] = 192;
               321 : lut_out[i] = 192;
               322 : lut_out[i] = 192;
               323 : lut_out[i] = 192;
               324 : lut_out[i] = 192;
               325 : lut_out[i] = 192;
               326 : lut_out[i] = 208;
               327 : lut_out[i] = 208;
               328 : lut_out[i] = 208;
               329 : lut_out[i] = 208;
               330 : lut_out[i] = 208;
               331 : lut_out[i] = 208;
               332 : lut_out[i] = 208;
               333 : lut_out[i] = 208;
               334 : lut_out[i] = 208;
               335 : lut_out[i] = 208;
               336 : lut_out[i] = 208;
               337 : lut_out[i] = 208;
               338 : lut_out[i] = 208;
               339 : lut_out[i] = 208;
               340 : lut_out[i] = 208;
               341 : lut_out[i] = 208;
               342 : lut_out[i] = 208;
               343 : lut_out[i] = 208;
               344 : lut_out[i] = 208;
               345 : lut_out[i] = 208;
               346 : lut_out[i] = 208;
               347 : lut_out[i] = 208;
               348 : lut_out[i] = 208;
               349 : lut_out[i] = 208;
               350 : lut_out[i] = 208;
               351 : lut_out[i] = 208;
               352 : lut_out[i] = 208;
               353 : lut_out[i] = 208;
               354 : lut_out[i] = 208;
               355 : lut_out[i] = 208;
               356 : lut_out[i] = 208;
               357 : lut_out[i] = 208;
               358 : lut_out[i] = 208;
               359 : lut_out[i] = 208;
               360 : lut_out[i] = 208;
               361 : lut_out[i] = 208;
               362 : lut_out[i] = 208;
               363 : lut_out[i] = 208;
               364 : lut_out[i] = 208;
               365 : lut_out[i] = 208;
               366 : lut_out[i] = 208;
               367 : lut_out[i] = 208;
               368 : lut_out[i] = 208;
               369 : lut_out[i] = 208;
               370 : lut_out[i] = 208;
               371 : lut_out[i] = 208;
               372 : lut_out[i] = 208;
               373 : lut_out[i] = 208;
               374 : lut_out[i] = 208;
               375 : lut_out[i] = 208;
               376 : lut_out[i] = 208;
               377 : lut_out[i] = 208;
               378 : lut_out[i] = 208;
               379 : lut_out[i] = 208;
               380 : lut_out[i] = 208;
               381 : lut_out[i] = 208;
               382 : lut_out[i] = 208;
               383 : lut_out[i] = 208;
               384 : lut_out[i] = 208;
               385 : lut_out[i] = 208;
               386 : lut_out[i] = 208;
               387 : lut_out[i] = 208;
               388 : lut_out[i] = 208;
               389 : lut_out[i] = 208;
               390 : lut_out[i] = 208;
               391 : lut_out[i] = 208;
               392 : lut_out[i] = 208;
               393 : lut_out[i] = 208;
               394 : lut_out[i] = 208;
               395 : lut_out[i] = 208;
               396 : lut_out[i] = 208;
               397 : lut_out[i] = 208;
               398 : lut_out[i] = 208;
               399 : lut_out[i] = 208;
               400 : lut_out[i] = 208;
               401 : lut_out[i] = 208;
               402 : lut_out[i] = 208;
               403 : lut_out[i] = 208;
               404 : lut_out[i] = 208;
               405 : lut_out[i] = 208;
               406 : lut_out[i] = 208;
               407 : lut_out[i] = 208;
               408 : lut_out[i] = 208;
               409 : lut_out[i] = 208;
               410 : lut_out[i] = 208;
               411 : lut_out[i] = 208;
               412 : lut_out[i] = 208;
               413 : lut_out[i] = 208;
               414 : lut_out[i] = 208;
               415 : lut_out[i] = 208;
               416 : lut_out[i] = 208;
               417 : lut_out[i] = 208;
               418 : lut_out[i] = 208;
               419 : lut_out[i] = 208;
               420 : lut_out[i] = 208;
               421 : lut_out[i] = 208;
               422 : lut_out[i] = 208;
               423 : lut_out[i] = 208;
               424 : lut_out[i] = 208;
               425 : lut_out[i] = 208;
               426 : lut_out[i] = 208;
               427 : lut_out[i] = 208;
               428 : lut_out[i] = 208;
               429 : lut_out[i] = 208;
               430 : lut_out[i] = 208;
               431 : lut_out[i] = 208;
               432 : lut_out[i] = 224;
               433 : lut_out[i] = 224;
               434 : lut_out[i] = 224;
               435 : lut_out[i] = 224;
               436 : lut_out[i] = 224;
               437 : lut_out[i] = 224;
               438 : lut_out[i] = 224;
               439 : lut_out[i] = 224;
               440 : lut_out[i] = 224;
               441 : lut_out[i] = 224;
               442 : lut_out[i] = 224;
               443 : lut_out[i] = 224;
               444 : lut_out[i] = 224;
               445 : lut_out[i] = 224;
               446 : lut_out[i] = 224;
               447 : lut_out[i] = 224;
               448 : lut_out[i] = 224;
               449 : lut_out[i] = 224;
               450 : lut_out[i] = 224;
               451 : lut_out[i] = 224;
               452 : lut_out[i] = 224;
               453 : lut_out[i] = 224;
               454 : lut_out[i] = 224;
               455 : lut_out[i] = 224;
               456 : lut_out[i] = 224;
               457 : lut_out[i] = 224;
               458 : lut_out[i] = 224;
               459 : lut_out[i] = 224;
               460 : lut_out[i] = 224;
               461 : lut_out[i] = 224;
               462 : lut_out[i] = 224;
               463 : lut_out[i] = 224;
               464 : lut_out[i] = 224;
               465 : lut_out[i] = 224;
               466 : lut_out[i] = 224;
               467 : lut_out[i] = 224;
               468 : lut_out[i] = 224;
               469 : lut_out[i] = 224;
               470 : lut_out[i] = 224;
               471 : lut_out[i] = 224;
               472 : lut_out[i] = 224;
               473 : lut_out[i] = 224;
               474 : lut_out[i] = 224;
               475 : lut_out[i] = 224;
               476 : lut_out[i] = 224;
               477 : lut_out[i] = 224;
               478 : lut_out[i] = 224;
               479 : lut_out[i] = 224;
               480 : lut_out[i] = 224;
               481 : lut_out[i] = 224;
               482 : lut_out[i] = 224;
               483 : lut_out[i] = 224;
               484 : lut_out[i] = 224;
               485 : lut_out[i] = 224;
               486 : lut_out[i] = 224;
               487 : lut_out[i] = 224;
               488 : lut_out[i] = 224;
               489 : lut_out[i] = 224;
               490 : lut_out[i] = 224;
               491 : lut_out[i] = 224;
               492 : lut_out[i] = 224;
               493 : lut_out[i] = 224;
               494 : lut_out[i] = 224;
               495 : lut_out[i] = 224;
               496 : lut_out[i] = 224;
               497 : lut_out[i] = 224;
               498 : lut_out[i] = 224;
               499 : lut_out[i] = 224;
               500 : lut_out[i] = 224;
               501 : lut_out[i] = 224;
               502 : lut_out[i] = 224;
               503 : lut_out[i] = 224;
               504 : lut_out[i] = 224;
               505 : lut_out[i] = 224;
               506 : lut_out[i] = 224;
               507 : lut_out[i] = 224;
               508 : lut_out[i] = 224;
               509 : lut_out[i] = 224;
               510 : lut_out[i] = 224;
               511 : lut_out[i] = 224;
               512 : lut_out[i] = 224;
               513 : lut_out[i] = 224;
               514 : lut_out[i] = 224;
               515 : lut_out[i] = 224;
               516 : lut_out[i] = 224;
               517 : lut_out[i] = 224;
               518 : lut_out[i] = 224;
               519 : lut_out[i] = 224;
               520 : lut_out[i] = 224;
               521 : lut_out[i] = 224;
               522 : lut_out[i] = 224;
               523 : lut_out[i] = 224;
               524 : lut_out[i] = 224;
               525 : lut_out[i] = 224;
               526 : lut_out[i] = 224;
               527 : lut_out[i] = 224;
               528 : lut_out[i] = 224;
               529 : lut_out[i] = 224;
               530 : lut_out[i] = 224;
               531 : lut_out[i] = 224;
               532 : lut_out[i] = 224;
               533 : lut_out[i] = 224;
               534 : lut_out[i] = 224;
               535 : lut_out[i] = 224;
               536 : lut_out[i] = 224;
               537 : lut_out[i] = 224;
               538 : lut_out[i] = 224;
               539 : lut_out[i] = 224;
               540 : lut_out[i] = 224;
               541 : lut_out[i] = 224;
               542 : lut_out[i] = 224;
               543 : lut_out[i] = 224;
               544 : lut_out[i] = 224;
               545 : lut_out[i] = 224;
               546 : lut_out[i] = 224;
               547 : lut_out[i] = 224;
               548 : lut_out[i] = 224;
               549 : lut_out[i] = 224;
               550 : lut_out[i] = 224;
               551 : lut_out[i] = 224;
               552 : lut_out[i] = 224;
               553 : lut_out[i] = 224;
               554 : lut_out[i] = 224;
               555 : lut_out[i] = 224;
               556 : lut_out[i] = 224;
               557 : lut_out[i] = 224;
               558 : lut_out[i] = 224;
               559 : lut_out[i] = 224;
               560 : lut_out[i] = 224;
               561 : lut_out[i] = 224;
               562 : lut_out[i] = 224;
               563 : lut_out[i] = 224;
               564 : lut_out[i] = 224;
               565 : lut_out[i] = 224;
               566 : lut_out[i] = 224;
               567 : lut_out[i] = 224;
               568 : lut_out[i] = 224;
               569 : lut_out[i] = 224;
               570 : lut_out[i] = 224;
               571 : lut_out[i] = 224;
               572 : lut_out[i] = 224;
               573 : lut_out[i] = 224;
               574 : lut_out[i] = 224;
               575 : lut_out[i] = 224;
               576 : lut_out[i] = 224;
               577 : lut_out[i] = 224;
               578 : lut_out[i] = 224;
               579 : lut_out[i] = 224;
               580 : lut_out[i] = 224;
               581 : lut_out[i] = 240;
               582 : lut_out[i] = 240;
               583 : lut_out[i] = 240;
               584 : lut_out[i] = 240;
               585 : lut_out[i] = 240;
               586 : lut_out[i] = 240;
               587 : lut_out[i] = 240;
               588 : lut_out[i] = 240;
               589 : lut_out[i] = 240;
               590 : lut_out[i] = 240;
               591 : lut_out[i] = 240;
               592 : lut_out[i] = 240;
               593 : lut_out[i] = 240;
               594 : lut_out[i] = 240;
               595 : lut_out[i] = 240;
               596 : lut_out[i] = 240;
               597 : lut_out[i] = 240;
               598 : lut_out[i] = 240;
               599 : lut_out[i] = 240;
               600 : lut_out[i] = 240;
               601 : lut_out[i] = 240;
               602 : lut_out[i] = 240;
               603 : lut_out[i] = 240;
               604 : lut_out[i] = 240;
               605 : lut_out[i] = 240;
               606 : lut_out[i] = 240;
               607 : lut_out[i] = 240;
               608 : lut_out[i] = 240;
               609 : lut_out[i] = 240;
               610 : lut_out[i] = 240;
               611 : lut_out[i] = 240;
               612 : lut_out[i] = 240;
               613 : lut_out[i] = 240;
               614 : lut_out[i] = 240;
               615 : lut_out[i] = 240;
               616 : lut_out[i] = 240;
               617 : lut_out[i] = 240;
               618 : lut_out[i] = 240;
               619 : lut_out[i] = 240;
               620 : lut_out[i] = 240;
               621 : lut_out[i] = 240;
               622 : lut_out[i] = 240;
               623 : lut_out[i] = 240;
               624 : lut_out[i] = 240;
               625 : lut_out[i] = 240;
               626 : lut_out[i] = 240;
               627 : lut_out[i] = 240;
               628 : lut_out[i] = 240;
               629 : lut_out[i] = 240;
               630 : lut_out[i] = 240;
               631 : lut_out[i] = 240;
               632 : lut_out[i] = 240;
               633 : lut_out[i] = 240;
               634 : lut_out[i] = 240;
               635 : lut_out[i] = 240;
               636 : lut_out[i] = 240;
               637 : lut_out[i] = 240;
               638 : lut_out[i] = 240;
               639 : lut_out[i] = 240;
               640 : lut_out[i] = 240;
               641 : lut_out[i] = 240;
               642 : lut_out[i] = 240;
               643 : lut_out[i] = 240;
               644 : lut_out[i] = 240;
               645 : lut_out[i] = 240;
               646 : lut_out[i] = 240;
               647 : lut_out[i] = 240;
               648 : lut_out[i] = 240;
               649 : lut_out[i] = 240;
               650 : lut_out[i] = 240;
               651 : lut_out[i] = 240;
               652 : lut_out[i] = 240;
               653 : lut_out[i] = 240;
               654 : lut_out[i] = 240;
               655 : lut_out[i] = 240;
               656 : lut_out[i] = 240;
               657 : lut_out[i] = 240;
               658 : lut_out[i] = 240;
               659 : lut_out[i] = 240;
               660 : lut_out[i] = 240;
               661 : lut_out[i] = 240;
               662 : lut_out[i] = 240;
               663 : lut_out[i] = 240;
               664 : lut_out[i] = 240;
               665 : lut_out[i] = 240;
               666 : lut_out[i] = 240;
               667 : lut_out[i] = 240;
               668 : lut_out[i] = 240;
               669 : lut_out[i] = 240;
               670 : lut_out[i] = 240;
               671 : lut_out[i] = 240;
               672 : lut_out[i] = 240;
               673 : lut_out[i] = 240;
               674 : lut_out[i] = 240;
               675 : lut_out[i] = 240;
               676 : lut_out[i] = 240;
               677 : lut_out[i] = 240;
               678 : lut_out[i] = 240;
               679 : lut_out[i] = 240;
               680 : lut_out[i] = 240;
               681 : lut_out[i] = 240;
               682 : lut_out[i] = 240;
               683 : lut_out[i] = 240;
               684 : lut_out[i] = 240;
               685 : lut_out[i] = 240;
               686 : lut_out[i] = 240;
               687 : lut_out[i] = 240;
               688 : lut_out[i] = 240;
               689 : lut_out[i] = 240;
               690 : lut_out[i] = 240;
               691 : lut_out[i] = 240;
               692 : lut_out[i] = 240;
               693 : lut_out[i] = 240;
               694 : lut_out[i] = 240;
               695 : lut_out[i] = 240;
               696 : lut_out[i] = 240;
               697 : lut_out[i] = 240;
               698 : lut_out[i] = 240;
               699 : lut_out[i] = 240;
               700 : lut_out[i] = 240;
               701 : lut_out[i] = 240;
               702 : lut_out[i] = 240;
               703 : lut_out[i] = 240;
               704 : lut_out[i] = 240;
               705 : lut_out[i] = 240;
               706 : lut_out[i] = 240;
               707 : lut_out[i] = 240;
               708 : lut_out[i] = 240;
               709 : lut_out[i] = 240;
               710 : lut_out[i] = 240;
               711 : lut_out[i] = 240;
               712 : lut_out[i] = 240;
               713 : lut_out[i] = 240;
               714 : lut_out[i] = 240;
               715 : lut_out[i] = 240;
               716 : lut_out[i] = 240;
               717 : lut_out[i] = 240;
               718 : lut_out[i] = 240;
               719 : lut_out[i] = 240;
               720 : lut_out[i] = 240;
               721 : lut_out[i] = 240;
               722 : lut_out[i] = 240;
               723 : lut_out[i] = 240;
               724 : lut_out[i] = 240;
               725 : lut_out[i] = 240;
               726 : lut_out[i] = 240;
               727 : lut_out[i] = 240;
               728 : lut_out[i] = 240;
               729 : lut_out[i] = 240;
               730 : lut_out[i] = 240;
               731 : lut_out[i] = 240;
               732 : lut_out[i] = 240;
               733 : lut_out[i] = 240;
               734 : lut_out[i] = 240;
               735 : lut_out[i] = 240;
               736 : lut_out[i] = 240;
               737 : lut_out[i] = 240;
               738 : lut_out[i] = 240;
               739 : lut_out[i] = 240;
               740 : lut_out[i] = 240;
               741 : lut_out[i] = 240;
               742 : lut_out[i] = 240;
               743 : lut_out[i] = 240;
               744 : lut_out[i] = 240;
               745 : lut_out[i] = 240;
               746 : lut_out[i] = 240;
               747 : lut_out[i] = 240;
               748 : lut_out[i] = 240;
               749 : lut_out[i] = 240;
               750 : lut_out[i] = 240;
               751 : lut_out[i] = 240;
               752 : lut_out[i] = 240;
               753 : lut_out[i] = 240;
               754 : lut_out[i] = 240;
               755 : lut_out[i] = 240;
               756 : lut_out[i] = 240;
               757 : lut_out[i] = 240;
               758 : lut_out[i] = 240;
               759 : lut_out[i] = 240;
               760 : lut_out[i] = 240;
               761 : lut_out[i] = 240;
               762 : lut_out[i] = 240;
               763 : lut_out[i] = 240;
               764 : lut_out[i] = 240;
               765 : lut_out[i] = 240;
               766 : lut_out[i] = 240;
               767 : lut_out[i] = 240;
               768 : lut_out[i] = 240;
               769 : lut_out[i] = 240;
               770 : lut_out[i] = 240;
               771 : lut_out[i] = 240;
               772 : lut_out[i] = 240;
               773 : lut_out[i] = 240;
               774 : lut_out[i] = 240;
               775 : lut_out[i] = 240;
               776 : lut_out[i] = 240;
               777 : lut_out[i] = 240;
               778 : lut_out[i] = 240;
               779 : lut_out[i] = 240;
               780 : lut_out[i] = 240;
               781 : lut_out[i] = 240;
               782 : lut_out[i] = 240;
               783 : lut_out[i] = 240;
               784 : lut_out[i] = 240;
               785 : lut_out[i] = 240;
               786 : lut_out[i] = 240;
               787 : lut_out[i] = 240;
               788 : lut_out[i] = 240;
               789 : lut_out[i] = 240;
               790 : lut_out[i] = 240;
               791 : lut_out[i] = 240;
               792 : lut_out[i] = 240;
               793 : lut_out[i] = 240;
               794 : lut_out[i] = 240;
               795 : lut_out[i] = 240;
               796 : lut_out[i] = 240;
               797 : lut_out[i] = 240;
               798 : lut_out[i] = 240;
               799 : lut_out[i] = 240;
               800 : lut_out[i] = 240;
               801 : lut_out[i] = 240;
               802 : lut_out[i] = 240;
               803 : lut_out[i] = 240;
               804 : lut_out[i] = 240;
               805 : lut_out[i] = 240;
               806 : lut_out[i] = 240;
               807 : lut_out[i] = 240;
               808 : lut_out[i] = 240;
               809 : lut_out[i] = 240;
               810 : lut_out[i] = 240;
               811 : lut_out[i] = 240;
               812 : lut_out[i] = 240;
               813 : lut_out[i] = 240;
               814 : lut_out[i] = 240;
               815 : lut_out[i] = 240;
               816 : lut_out[i] = 240;
               817 : lut_out[i] = 240;
               818 : lut_out[i] = 240;
               819 : lut_out[i] = 240;
               820 : lut_out[i] = 240;
               821 : lut_out[i] = 240;
               822 : lut_out[i] = 240;
               823 : lut_out[i] = 240;
               824 : lut_out[i] = 240;
               825 : lut_out[i] = 240;
               826 : lut_out[i] = 240;
               827 : lut_out[i] = 240;
               828 : lut_out[i] = 240;
               829 : lut_out[i] = 240;
               830 : lut_out[i] = 240;
               831 : lut_out[i] = 240;
               832 : lut_out[i] = 240;
               833 : lut_out[i] = 240;
               834 : lut_out[i] = 240;
               835 : lut_out[i] = 240;
               836 : lut_out[i] = 240;
               837 : lut_out[i] = 240;
               838 : lut_out[i] = 240;
               839 : lut_out[i] = 240;
               840 : lut_out[i] = 240;
               841 : lut_out[i] = 240;
               842 : lut_out[i] = 240;
               843 : lut_out[i] = 240;
               844 : lut_out[i] = 240;
               845 : lut_out[i] = 240;
               846 : lut_out[i] = 240;
               847 : lut_out[i] = 240;
               848 : lut_out[i] = 240;
               849 : lut_out[i] = 240;
               850 : lut_out[i] = 240;
               851 : lut_out[i] = 240;
               852 : lut_out[i] = 240;
               853 : lut_out[i] = 240;
               854 : lut_out[i] = 240;
               855 : lut_out[i] = 240;
               856 : lut_out[i] = 240;
               857 : lut_out[i] = 240;
               858 : lut_out[i] = 240;
               859 : lut_out[i] = 240;
               860 : lut_out[i] = 240;
               861 : lut_out[i] = 240;
               862 : lut_out[i] = 240;
               863 : lut_out[i] = 240;
               864 : lut_out[i] = 240;
               865 : lut_out[i] = 240;
               866 : lut_out[i] = 240;
               867 : lut_out[i] = 240;
               868 : lut_out[i] = 240;
               869 : lut_out[i] = 240;
               870 : lut_out[i] = 240;
               871 : lut_out[i] = 240;
               872 : lut_out[i] = 240;
               873 : lut_out[i] = 240;
               874 : lut_out[i] = 240;
               875 : lut_out[i] = 240;
               876 : lut_out[i] = 240;
               877 : lut_out[i] = 240;
               878 : lut_out[i] = 240;
               879 : lut_out[i] = 240;
               default: lut_out[i] = 0;
            endcase
         end
      end
   end
   
endmodule
